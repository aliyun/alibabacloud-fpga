`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
oBXvm/W5ec1IhJYI0f+5YaboHfdb30es3D5qM1mIhJ29UYtRUqL437Xvqk5SsidBjn8Ls0hMboI3
xRDd9Z/z0w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Hx+4+jZ+Lv0Zv8Edm/ZmizJ59xDfFW3dZeSmJ0YUJEDcYTX53J1GvWzXX04aYHWNognzNFFRq0eC
JTbYFGlf8k+LZRnyEYJA6eOOib22OrBbMxbhf65gQIgMOFVFc9SXOFd/cy81PIJkZ8gDRIMR5gAL
yLP4CqpuPsEnyBrwf+0=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dRq/j1bLujCvSMlBmMnQFGwC/tSWXEWgu5bvnI0LJt8G1/yFAcieyAquhx+n2KrNFJAwUtfgj0hO
jzb3XVpwy+XxSj9og5mwsohHA3/dWNWrsBpuXlTpvVGprxBWulLsR7+SkLBKLa5lK1C5M1kaa0IE
/GntNnn4a6hYHYlXkuEqKn9dypDfsy/Oq9B05cdFiUqr+vtvfySimdDUNl54RHXc3Ot6AImulOAC
e4pC5dwp02EZnk/2aUxDlDeB0BRRePFUs27E8khAUNRRBc+POYVpvLJAElPIr1FYG41lejMwz0+h
MaxQ+KjYobicS+04CodUIPFFHyocCCc431klkg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vN40CR2WDYkFImOzeLoVAlDN15J0LtBfAnMObXH6Bg8E/f/ZMSjGorsnpNWapJ0iF0iTS9BncSiq
bo0rHjJi1D4w8um5XOL0G511PIo1hAvYzBA+u+5WjjX669xkjUaKuZ2AN9mthC8xGTl3EE6x5rhP
0cn8+Y09CzFlYIDIOlxrC6Vhn4991CWl8jtpBMZ6wQ7LSnCOG5YkYO4OBuYDrrsaDMnvPmqhKv7M
ymRJrW51zKG8GqUSUMu99M/GQM78jF+ajhBN7iNFF4dM7bBW9b7qJDyrsQwdAbORrumdfRX3QcpH
UX5zeC+uWQk2kl1uoc5ICNPx80++RVXtPAxspQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dO6WGdxAulR9iqDJ+Q5xAthzj+Po2qkHp74nNiDdfqnL3DhKv2yFVv6zq0bBYmVHjGfAMJf8+uHK
rKx+tW8p6OhyC9hGCc9Z7QbjE6iox/i9vG5Pp3NBjR2uaLmcy0w787OmIYqAg/Spf7bByccBBq7i
nNt464gVQFlAUgVXHq7wYkgqdH6AIabCbYuMgiqJ6NShpcGttTsKp8gC/q7bi3sZeJFyYzeuUova
+Y5IAfGs7TvcqJM9BalsT1Aa1vTMJUHRYYOkcusNcyeAkLMcRIWQn8pPT0o60m3yrbJ0fm6VDQFr
++8lPAitCLDfGwUEqYfek8obBHTpPYMDy3xAQA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
rULiW37wBNsdCsspJ1o7aYGLHNbsnaKHpb5n4PgfYis6prtTTWyoYmQrdP45ZNLQNCpEuPOjpeqO
hpTwYJY4JIort/H/7OJTu9QuAHlu35CiI3QQxRM3vFkG0iVba5ZSdpcd1bU1TSrJociY3SDmajQg
5xP9f/JDgHXmMl40Ods=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MZkItI8j/BN1sxQAqBxRTKmPCnoOL2MmS6e+IaHGEuAJPzaKXEvgjm2/GUnC0iXucYViC4/BEW6D
dUaDqNv68zfIMkBpi9i7UT78xv2Kvp8AByCqsnoSDM855KdHSS/Q9UCazOMXuto4fJUKNqvsJaoY
6U5sClWBzK7LF95JMudZUciwmMX1WjeWt0mNSh8luJJ3ku78NW/lF55LxHjM7+tKPQ8LPcvcPwJ4
quL0+KmFTs2vcwAsIFRCG5SVAAcRqYMMsEYrfGP47nC5nD0BAy3YySP+ACwiGDb8ZPTMb4l+VKVP
PGLQwS0mjMQ5DBKCAXxKhKvjJy47LlWEv5UAeA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135968)
`pragma protect data_block
1+cOdCWvhsX5cR6jlD6OilbvY4SI8ROc8XcLh/NB/i3zHkez6j5mGWS6HdKxzx0apM3mu7ophAsY
o0C3V8LQdLseyujg7GyPcgXg+V5PzBFP8n8b8VVWQZb679a1vPAbDmSkqdpbQ9XvfJUBhrv0ipQQ
papk7b+SBIJNejv9WRKgtjv6ZAWrOhYweyIgysRvHOVdJnHUWZYwtUsahVz9fOzagQ1alEHK8bU+
jlkplurXQgEKy2Kr6dAnFYiCkgMgU/hPzaa5wmTxx/hD4QooGJ7sH/hWFY9wcD2xOaqSNzDBIkDo
AyPp5vVIFc13wScFgRP1Nr962n4UAlL6G1pcW778tKD6hJot2K9MftGTYMVM9ViZ+1qYqhxxouPf
ipdpwfq7wpVg/nuHsU25vMpFShWeqjCfS+FzG5QSqz1Ux632CZ/AWZQL979/TSV3DptdbDeKIuKC
KzdyrCMa5bAA+SOPzfBTm/eO3m2cexpaNRyTvXLvOKQbpg93JSFuEyGsJrJA1XyJEXBkOE4KuJ+x
JJ1FbD/WH+1QECu2fG3rNmjW4jw9M/gW8uXHSFbluJzzUaL0+Pt0GLUxbH0XPhQ+Ob3XX0WCf1n8
Uhw71+puVgYrGIn/BCJeDg3WU6XYKQRguMmwvB1AnYBI+XhH/BVy5ktCzQNAVrdcd6RX+rlxrLri
jHColxdwNi23NuGFcgEoDIIDpjpac6dCggmZgTra6jOrrt0BERa3TL+1c3mbLTK3qUNED3UkGz80
mIPQdij2lrwdubvQIH7Xw0L2OnQE2ss0b6zwOkpqeZIH/S75aPWP2UIKzLpigdNYOl0aCjOrC/vx
23tTlhuc1jjDJHk64+a5sppaT7tnIZfJ/Zn37WEKr59bVD4iWJ9l/yhMFAUy+hilIeMDG032PTRS
Y1YasO7zX3l+G4ChGx3yT8lMNT8KUX+SGn677/ckRmOdvfNY2PedPZJxQZrvgHuUxjZQDWCnhcIF
lcyjFhZ+15WAnegxv5qFEzixT5U5nsD142+v0tAX5T9tOWqwAR8TiXHuU2qLaR+qt2gHELpr/g7J
w6ntPNsvobx+pQnd5q3ZmRBX9Mg3r0NEZdBKx/CGeNiorU5WkB+xcYbLxl3OH8BRpyswn+3ua2UK
YJ49/Fqn9/ROsWl9g7CqQTPxSlRU9wxD5bAQe/HmGVXLEGsdF0zGsADO4GjAJhnK/9N5Xj/8jsKk
fFDQBVkl/OU2JBrH4TBdLawai/ksx0gWPr/NMbXuOGCPkjAeF++5YIpvH3woqPMjEffELYSe/1+q
ca3AYvGmyo3rZVtFwKyOpve2QtbxXZS6AumF9mAm8DuN3dNSmS0eWPEYvCfU7GuPTLFUTJAA+isk
DfkI10XTWSUKOa/xfEvGfBt3p5tponlmWppoHxfEpTRXX9o95gsZWGrmCcJ4xFKImB1hfjz1ODCh
VUBJ7qBDO6FGimQ9bBwxbJpvAYaFvbUmjEn1PQ9Bzu7X6KcAnfNQvrX+ZFp1l204r9NlTQtMftXm
+TzOOE62lJ/gspurFn0jm4Iq+fbghb5e04NUiIDCwwgAAr4r/wtjftGJJWsJuBRZoAb5kT2JdSA7
4qInFnqTgsOKQMPER3E7CgJWwzG/bXEJQAfEbwz/WwOkFNBLwwjPC755DA72NCrpiNpGZ1LeNiwZ
zVt5FSCexaN6uwEuf8/I0dCn5f7614zoQi5YDQuG2HgfjMDdcKF4yipFLQJDSep3e/Z43GXg75bA
B6p0es+yI+EhlOVw12pnz1DrWc1CR7iXHkJ3SZufuorRIob5NgEv3Qw1cv8gvWJ+h2k1BNVRU6NV
MUwOgnVJCij7kwtJNdkIybT1hs87lRXotYiAvkUlHZOQoR+L5VUa7wegrfieesan4oZJqXig/epo
0QsDpMOfdotNtGuaAxZQWaoBwIBjeQLXRpCJY+pKcXLgseZOCSdxlXXv1BOv9OLC5eJTTjf25lsz
jwX3MQkTNEA/0O/9VXxmmmwEtpgEa3fn1Ul5Hco0HarGGGyBbNG04cvu3iEj3wI563i/aihdfZUj
+lI7hz0X11R5gDhxMwrGy0eTe/BleX8UoA3FZCWQ4gbvESbzE5rsh8NaYt9W+stv/J74tR1qLI2e
LzQks2Gk1h/lZG7EoTEkIvRGkAbwbHRUD6elnheV/tpI/aZ8yvKWuUotWuCXhRm9emQcz0xZ8vcS
uVGSM86qhiuBmBdenBXcPbrnet0FBZJhTxo70CRnDIkQxC2uLrpn5OZYi69iMmSx9YP0ptDGBI7P
t11rUILiaxJ1I2gk9PS3Ft5MJsr79NbtKXGvIwkJ5RWsXdFjVdQAXelk0ANi3NZOafU3GxnlNxxn
U7MbnaJggjl6zyiQQUJQP/8SaVI/68NYsTZ5ZBMhfugZ7TpfqYSxU2YXQke+XFNTOKtlM57qFo8b
z8EauirkBX6Bc54UrP7aktzxiFqKacQPoJf7ucLoC7lm4PKd9D/D0WFxtn9oX6EmvUlkmSAObO+t
qce1d5YleQ4+/yEe1d6V09Svqo0G1lp9YJExA1JoS/h+SvS+eFUOY1WdQP6NH+OFPgLCbkAkMxtp
U8VwUyv2BSGAio0iKrCtglb7wbARLgrBzRvtGyLPzWr/gGzbjBUYGHLIJZIyuAlZndq9/JXn+Osu
6O0vagb1Go0Fx/h+fNYtBF6xtMCsC/b/+xdiaHK35ssfIHtxFgHrJ4Z1FO53grYxT/26EIdMO8Hl
F/GVGcOr+aWsvs5RHl1S4cOzueq+PkpjEL8Skvk9mxJ3paL4y4H3DbD1rYUhzOgF++rWdVG+jZhL
2aI/VS2RfZ3PcaDjolj8enhPMg+Kfk/L3ykeqVvbpyP5uCWYBGGTJXYPwsmq6rHDR2gmez3XIK6K
nmoAEcqvqHu5054Cl63VEH2MmqPjYUZPq+Y08HFKQPHYuYCja0mbk8lESoHEQvx0b7903OhjWBI+
ZpjxVMT9lwSuLaGrUZmiLwNc1VAQIqQe70EyiOyNOgROCRj8ght0uS60qhSH3EgRnB5LYRs/kKai
uAQA9L/POUNAlKZOBA9ofv75uCKEAB9nty5u0r59uakCw50qUHzsT035ztQDILzUKFM0qXh8c6oy
FkV/CguAA7a5JFtYwHtP2vNuq/5BUUxvvr8mUIozCJ3d+To766Og9KZ+wLMhe3U2LtTb+7CewmQ8
MAZPWdyZRHL1sMxV7W/CG69GQ7thW9RmplPq75I+iII3DsefGabUCM7uKREsTRmvFXIyWSzvSfmO
M4BUB1OPqFxvB54kP0TZG8qTjRnG8zgvv8bM+vCu7165OavV302GUc/gBW5eLgyYRUbC7NZN05eF
9v/Slx/JVUNE2FcazOhfDZ+Qn1XEXQqBpSPHy41KyOwu2m3AcWFh6acTRa+we6cV4qSSciI2pKqb
JtKpzjWPd2im7FmkMSCjoIs0B+OO63+xn2RBHVAWTTEx7ZhiJ+r/N3WmypqybAXEnzayvut4jwa8
iVUTu3Npz9NnuSiGZgT0+UXjW7j+xOtyli6AnjOqNMTS0Qe8aZ8ZfMcBSMeOVFRud4778c4QT40f
Hz4jVTiFXbfY/HVRwz4lzgoR+StXumr1vIHgjW0PW9/a6hw2An93rcslS7kIWzkk/enE3DqReWr7
vXDFTXygFjflFNipPStLmA6wyiYxh60zS/39jz3gIzRSjAtIq0/9iOsZw8pzxAdKn5ejXkdRQ4s/
jOgZOgXOQyUNn0O2JAY8iV/VdqyP0MXic0h62WGP/OqLrAdVsRgnrn2vjfvuHLp/JOl/ERHa2lDJ
2jOL0ZgUGjCeSMFIWgqcbMzTcif2s8ZylTx0IhvTJLXQpMlwRaxsMImH0CojH8+qhSmr/ynSkDbL
uEbMH6gXsbV6u/WC7LVulPGPW8PIH0+vIzZ7omGzRm10sGy/gmfnyAoYw7OaaXLURGsW055v6jZ0
O3iqIjM2VPo09e4aDqSGjdN9uuXsKabPhkneYBY48eNsYEb6agyELK4a94i/9rO3I+UUqRRuirVU
ue6F84dccNZ8hTOK8aaYYmJx/5haptbDmFtO5VSymgNrCJhAvEgAyT9KxyXL7r5tV7z7gVQHlvZ1
ERHFiZyfV90WKGKjpRIBSy42TxCnjt7KmlmcJYpvzwP0eWJVNPSIM9C+z7c8iOQQU4DABxJXdhNo
GN3NEgHCqcbMO/4AGNMvyVSrmoGqFXZPry+kBu8Mj00lAzCsmKupouleJAbALsjIZIiy+EsKDQ31
/4BrO+vwLb5SOcJxkIZIYvLi09Z1ktGdEl6FsacW3+7jgk6ICMbRwz+ykzYKeAZqVnePrybSDoFM
gtqXNN0i4Fq//Bi9zt8VYdP+8Schag4cbdxMv/FIxjSd+eyetkQuoP4nxM3niT6S7VjVJKPpeuG7
xu0HRcU5LjvYxauVuzeGzAlE5cjTKxSfTVANZtX8kUGcQzx6oH4wDjd1s/JoWluIZxMFMtDXTjjT
9fwn7w1KniJyF6mFo1hwsJ2PssOQejfuAEaHY58BFGvQ1Blh060m0d5vqMYWYp/hrJxIyvd/9kXO
UAK8H1riIhBCLkTU1srmRcABQkWQCLgLTIWEZ9Mqc8TCNcZsISJuuh3E2RIzwNCxQu3gQSE1GRb/
LMcmIRiWnIA4GgRmYL5K0dRsTXV018Im+xnPPd/K/EJ5VrvgUGtmrxxXQ8ax+onTACb38fX2nl8a
fTjvbtyuHjr/ei8xRpL+jGdpqcdrN36WIo+4CC6SX5RYqB2kMD/sQ3vuDjx+jjEydXa7hXwzvkJe
U9FQX0cAEFPEFjMBWeAmh8hbLjXWb2nvj9nfPfSzwzeG/YqFzbM+TrvRKkXRbLSpFvHg4ccQcScz
5f0N4OPpMB5Bi9qViPE71GkeMQOil3VxzGEYXQbaPm5+aD1jg2zUhA9krujfRiuzS44NO6Vb5Sfo
LWZ/alpQ+tSXo9MLLGMYusdk/kRAZYNV6DSqrTDiXaS6XBVzvroW/2K1pUVj2HpAVCcj2L1dAXkj
sjHv6IKeabpTvhKzAx1EYsB9paSWnBexb7/hT/b/vQ+P9/72X2mepB113GtoQCpoGUmrT6onDrj0
7as/ihP0LTJZX4hh4/A4d1xQPkWThwJuyhdY4JZbbkqqPx4DDiLcloTPUP5Lej58vFTQQLxgNmtL
nko3UsrDiuEIXWIlOJmUOKkioCT+1ls0Ld+S3U99GsU3EAoZd0O74jZE9LVxNSa+4SqkDoN1OTVZ
YLBg2a2ZNUKXYw55P+XKCD8hIp+QwUizQJXb3qVaVqHkvCWA3SsRA6JEdD9cYhln6ji1eDOyu/9C
BECsGQg+rSd9l5hIqg30Gb8/lYVq9k9PSYYgVni/pwLXu2oYvB8a2HLXSXZw3IFAEYLo1gJP1ScI
nP1mB4T8XzLsNBQCRJpBLM6emTCmXn/gmGl0eUt8uPKo/x83+qGjcFS96lpbg2NlFVG2Z7W5/1Wf
P8orv9ffZXx6Ad7L220GsNwZdZyq8ReSPJG5Ue5O5fJxxl2hDUF9ljNMxK1DpVJlJQdDnCJiSqhj
UnLWiRubk4w2vJGXP/nKs/fT5WEwmu/4TDhL+5g1mFzgxp04ff1nFThkql+kvHwrbAtvmxGUzl1e
FWQxO0FhD25mN4aNU4uIQ/J5GGgtmEp0jthriaPjLrThyrPWjF94DmsOkuCR3OkmI7pbZBnn8lNX
CSXH7/TrXJ2CzIS3XfT9in1G9fP/VL2MvxPRU45UOFQ0VLj6uQpcBGvxzB9IH47tDWv8/trtEmg3
bUafkEqQtDXhMeopgHubkyt4kMdV32e3z5B8fd0vidEG6ZOsHyjOjXnjFeQQAqMUT9S9K7EU168y
+6ApU+kMi3s89C8H5Gn8snUqaTR+Y/HdRIiZeLdGXnSdkHjt32oq7JBjpkCFAUYtfdJeaWkqm3UU
0CYn62xh6kCzU0CPk1Mnb1qkTropoWIsRpENTXQbdRDCOR+J3OCqDep9ohHTHIH6OJ4vpciIdh1I
/wbQReXky3GM9yokBJcGJaTPiLthTrDQfJkP5pY8ZY89UbeXYDBQ7n3beB72HEDG685aL6I9xAGh
oz1deBzuFW20r40e7H8WWxqTXm9FpZlvhLOfJ0ljQJIcluE/0woQwhASMoKg53nMG27bgZvys20c
RuPXjHXzT1C5z1AVpv1d9LA779Z/5zHYnN/A5nhEev1rxap7JeGN6wQv4Rapovf8vgyljyIxHr+y
6gvSFGXlWdGIDisodvobkqgIeeihbhpt9Z6bhUnG3bV1j0E3PvbDNUdKWm7NblvzMBpMyCFE2li0
dIpBJ4F58rJn5VxDulSYxzDbnNWAFFVZh3MC6atx6/ODHLtJQLPY9jqEJvlFSfltr+uLjdlNPPZh
jNwD7X/JHRHPTrTc4TMX6M8Z1MjsJfavF5M8TzcaZT6wUhAvUikqVOIeYGw8F2ib6zupbDiEr2as
i3NfZf+3eIcKQPfJjUxxJyoIaJUKAYCy6/2PE0rohHKRVJKU8QPO5gUtGlNqYkUArATCXclIWLyE
L96Urps8mauWb+TdNM+eVDDL5mrfUTwxcBHemVXofRRrd3bAlM9wvl/dm1pp63evXvVqIUzoDO/2
9ji8l+tCXvhHdYbkoMcx6lafhaUlNq0O9+5KbSAf6dtRD8db00wj3WVNwyk1xAFHckS3PdHLfkKZ
B4TGx20RrGadBGQTBBnV9bDPs8YAYqwf3Isj5Io+0b62ORp/D7bnC62oM/UY0Z0XHlyoOlmHibRS
sSWpP2QmXPu4SulQaG8r5bcvgUL3HbGAAGm/Y5ipmKPCB/ErDP+yHMvEkNsuXBiN4yL+/HZeik5y
VnRqj80o8eSC5WA87LWYlchbF8JucT131S7akXcZh9xMWAgyz51Uk0SwgzcMGtHX6Y8KTYujvuSI
eTuYX8a0srJKIUdj0lunW2q41HsnlEKPWuaMzrWM8A10mLL4HfnA7aXvBs6RRCP3/Svs7LHxBhBc
OuuVQYDTHXdgXfmyXfGVOjnaF4yPFOJA8/13sBPHJrsF4lKeL2dQDAUo1yWFB0bqSqP8sjsl6hBN
sd/UD4yHCFM+Q7IkV0YOUwYXdrAVxCXkbEybd8VkUnQDcm9bdNmOrOunvxpxlMmN8Uhrgk2MZgQV
74HsF7KEX8Hm8wvMdfcVzSE8qZkUmkfDR1xHSuNGgN+iclc9HLEuBIRzLSDb09iZRa+YFb9zMD4y
85oFOI8/vUbKpsLDVH/J0nEnfv6GNc+mE4zj3KX98fkA+LfKHwKyblS8ibXqjOpElVUXvY6EJFyH
fCU61vQtdmUg2CBUyQtfgkAvNghZqfwz/GPbuQQzlujy47CYfewvD15vfrNyQ4ImeqV1/6y3mmnd
tNTvQx7Un5PkdomhRESKcRslEoHDcVwVMiyZMwWbOvrkiL5Hsw3/Vzy47B6IwRSxOB0tQBpebows
L+LRRqOiUBDlWQu/INtuk7UzU0qxKb2+qOWZHyuQBozcuYTI2iyHrna+jVlw7/qQwG3eYjBfuJZe
dD6K9QWWSeCnVMwtt0WAq+rbKuuMFrpZmPHP4Ryfv7AKKu3uOwAAFBT12m7uhyvYatCXu3e2vvri
bsGswD/B2FLCU52XT0QLHrYREbtUuIjO+RTWt8uV4hzIfeHMI7J8AaYtBtD5p+yQLI99NFqEUa8/
bmhZKu7oxF+fSol/wUfsTgh14vK1KN5tjZ6gpiIHjaxEOvP0WhFyM96zED+WEClLPYkui/3kIr6f
Q3CasXHgjPDB30MOBSrY+vSCHTGEW3sIRSUXuOMXnCbN/MbtT2ZdVrm/rgo2wdadP1LD4SZDTRc7
aFdYoeqBHWixT5tgwplua+RoTs2sKaUlK5Lz02Fnr1VEkLCo1e8Dsdy4KpyS+7nNYcyqIEbc6Fv9
cJxQejWVvYj7/hz8VkOCI74pa12wip0IEN64RC7SppUwB7zOwpqqV66o51gf9/g2eKyFqsi+MgBp
tzL9GsBZWs8RQCTaO/hmzWeVkZnMiEkEmV7f2jbNhFJS05spTARCXKyIttg6xQpyqjHZZrXqdmHD
oD5SqXIKf2FthCs1VGteHrfa3wYiauzWI3dKxJiO3gjjRuWvG/6iCwm+ucqy+flVZC0sYoNk/SmB
uZn3BnYbSuQs/VqU6kz4dSKJdtnkXCHLpZLTAbIPHxZYoY5085gGpLT878Q4CdUgG1cJBiqDA7fV
bYuUuunjZW+ICO8gTrY+q+5ppZsRaPGvZy9GilZexGpKIuC1CDtuGVu4Tcvbx0Q+1QyhjxBZfpl3
Bwwg/pD9L/X72FL5Giu7w5YHEGhgzJAh6wkATCpnrzQwgPJf/lRb3rEONRUkb54NIf1CX05vEsgo
QUwBpfjvnbNQaUvJgfuubjTwoPqsn0H7eDvAFwiTmGMTKq4jfexopalFapWYTLyPAWdkgc5iehll
ibn6zjjHDYhjq6EMhpC8r1mNRFZS9dp8AM+naYIgCKsmRcGBeUNgEwz6AJbcU11G3QYD+jsOtb8w
O/1YJtw0JkUQuJmYgJbtfquNW+bM6iECEUNNBpS4khQFuB8D04v/pyCkaa0i0p8DHMTQoq0aNgLX
SETdWewqE2poamWbomPEBnHRmRPEXJTio2yWKd1nKwmRWnqEvtWdu9spOim0y/ZHHhKy/aRzdvGW
bFm6BskDDjLBUkTQc3M7gshYP2tedH7W2BGiAKH7HyQnbl2/1Q9gRYHnRXqBiVogqqC19ebEFqgd
DvT5pq1dNZ+/NcUAoprWQVBOTAoiHNuChKgl7bYHITxDG2p4Y2DPaM7ncH+hXNg9Q29Up6ikXSUD
L5BXWy5Vdeux8fQXnbiNedFZXc5LhHxy2PF0H+N2IBoRGpbeacH8+XCbLKIAV4d3ZfOgSviA8g3h
o52q2OXywDW4a+YU7XF/lAGUEEBg9uUOZCeGw3JbWXDdE8x17qJzXNsXWuiNI6JLRj17qYpES39O
sjlFIsaXEGbuP6PRCSxVBgIUHqJgYpHxnsjGAwQhPF5ViTNPXxcnbnRnULNPt2jeRnPrhFNLzIrZ
Rma114xU5ShO5L/OG4cjvYwxo9SApGVHMGeEPh/lt6C5Hq1Zoh2gpbtVFUTpQOz52KHod99nbrzG
Ryc6Bf081oaRCbULqnJ3zu2Q7Ty7K/kFHZ2VRu7y5MwZGd2Gw3F7cjHo5dy4sDSO+bttjcR/sWwr
cjKzbzXS/0f6FV1L5g9fI9HIjLjGEnT4AmSfVp0Ln4Njn4vO6DJCAxIZer5N+Q4KNoHXLoXUV2xz
PwCswlrBpQBC0Fd4WE/CMirfxQGkgDd4raos5xskiT2vd0Ed7vRAM8oLzQ5b2SdxUnYuoledrLwH
76fbIXkxkUEOecCxST3Tw+YBG3ttCiougEfAuohXqZ4GBAJ3/Hv1u7O097HDiNB++fAqNBE6t7l8
ubI7qrivgwasPUlb1oVmyB8FHfzsZPg3XVxrZNWe2R79+LZB8roUstHCUwQDkNzTRGspr+s1R7eN
SHyxUGxYCmKfBlBpsFarvyoPCmMXll64EtZ/a0oC81dUrLaR1B6/YYF136qgm6nw+CwpkO0N112n
Be0OfJ988yy7BFHHqQR8qYvBDIm4cqYcRujWfejW+44vtZZBp3HrWkr8QJ6ucATJJAElJzN0DpxR
uFChSE5XBTQs5ZvWoWDQv3uMIdRBE/xkv2kEoOvsSjuVlojTPIwbWfQqxypgv7JoccRQhX+bYqB2
dS/mrm7zPpv/gZGmRXn10v8nCJhtgqTmYLZscHxc+RU22ITgDonchZL/yL+47hHmWbUrxg3Ekdlk
OC/MK9j0W/z7PQ8cWQfXSYr1MYXj6jZiZ42G6WAclU+7hETkkUmcI+h9MD2xTudX9tIy8XLCDuab
L8aZSNgIMgb7MqEFFnygJp+Ym+iv5An/vgaNJCcLUeMK6N/ZkY5sdlXzPgQj7x1jAMpuW+S70WoU
78ChLj0aejU8pp2JfIhJD6kz4rjJJi5R0Df9Id9Mb8ZYxpBnzfNPOhlsDScJ4BhrzIGY7lsKoyyw
lP/3cfzjVta0VhyZ0dYK2Y37TAyhZpETkLLAOPKCpehuQMvJV6EvC1KsqkfvcQKNYOiMcYhWd4kD
FYPdLnBSYofnV1qms6U7zxvbvU7uH80UbXrJ+4gRZYBqbZvCT0Z3Q79HGaGotxeEfcxdG1v0JCZX
SsLn6Wciv6AP503HQf/aNoJB6vxcWGg70+C4ds0ySOZsj05j6TjS8HWe0Hm28qHG4nSGmSC9c/5q
8pWWDPrIKVmxT98+90RcuLk2aWRLJnOdgwX1EsbASNxdRBa/ibZsJAmrep2+SOCwNbArem0RJtGN
/qv+K5MvimgeX68ZJu1SbGQp3UShkn/NY8dzZc0t9rcBE6kZ3YqYTR5Dg0/60y5ED+qb+eN1rF+4
k+objQho7fT5rT7Awgaryhj54NFyHUtvumV071osZwwzqJHmBn1Es+psV7+tvo3yu0EFrLLHXBUt
fxE8XfvpKNfWpnC1FvoYIiSX7PSA2lpYlx0ZtnS+bOwmFPKUVVr5y57FCiM405uRL/5nrrMbV/Vu
DapfS7HpeyBFqIy3sdlQ+nOq1mR8CwpjcWFX954E7d+m/m+/5uIKhNBmDH+DMk6R8UkhD8rj4dmL
rz3ZuVSBfsBsOrL3u+psxU9CvfJIA63vsC+I33ygJivel0/j4SGLnilR3iIwPXJ0zvSt9slj/wpH
OXC1BX9vPXRgiCaRuBOSS7YWhuv/mcK+T7wEEyIM/VVyv1zgr7t00lGJycB/8ufTDoCEPr4Iyk2U
LXKBB1pNv5/9aZziWsSoiO5ipNxBLg7JdhHXDjzQIgLV3wFHcpnajBkLxSkqAWXfQwoBTk3eZ13h
hCSE1TkpSFmgPFYCAfLl7apnV3zW1RJphcV1Zmi/h2IcqOUvWG5l0yxPOEfX0dreWvsNE8epflte
5y7LFt/rZwegjgjjad2kheAQmXO9hhFAERRUAKNUd/1ihohpigyR50DI1aHrTUpYs6XEyIrRDwL2
W26LokhWOMxvkLxLS/62J9AIaO6dqFo4VgtM359whZZN2F1LCIrOPdoKPPnmp4nnH8N9DWMlxghJ
3IJlqakEd2ieu20jpAm59SEN54aftE0lMD8vQ9MjE+iZ9eGknYhoQkkaflw9lZtSlkZ6T40u0gnc
4czodQQC4BkCPVyq0Uv3WH5WatSTBQuCrOMMFRoGn2oGayZGsLBgHNp1BVk5A9ipOc808a6aaQEp
59ElhnH5Mjudp6WXwxIKhLG4a1bMuOSHQDZhpDkLS9q/oeD3QRQMmAWsj4nzUJRZbI4FvCSkRBwz
+E6n8UuDZaCL253hm9IgaGykT01Eti038jocRls6puz4B5G/wbeQIsMGVW9j9hu+4nADlsYE62nn
Sk1FXf0KCcP72KY/yRQQVxbQU/AEHEUqCHL4Jfq+JPpI/BzC5Pgo0FuQk4kaFoAw3WHO7LxCMIPu
uUzEko7Z3HWVwvF2hvRWsk0F/jEP/eM2HzFECHs5A4zYd/c51kiJFDr1zUKXjDDOvI+W81TPeXk3
L1SJKfjeEHNgZe1oHHqwOWKDbSZnSY30ddHdCKLtBd+XZUUTkIpXthcoPAl5zkz41l3Fv4YvmJnP
FwaF8EHB13t7DkfjJTIxsA/dB+wR3FY8EHolAvRjuR285tCU2FVmEn0cgtWcd0oe6CrAKF+SmEwI
tnAQ/jQJulnW0Gd8dMp//j2XKAaug06MIMcrYLNTLwpYQq4c7qcZvcF2pyP5qFY9v1M559DFfQ+E
+L/SguLyhfnTjaZV9AXEr4w/m83cLcKB/pNb2UdvU8bEskss3Fd0ECKRIS9ZrenWqGsMB5vI/2se
hLDhuhDKuDGmu8Q5yFtJtmRWh149Mq5RAJb7drRpKUD099YNUKFEbqJFZU+bOLb5K+pD7OzyhCh8
vYOTJpf+8GSkmmIieKmzURpHtmk+sSXiP4o+nFzuzJntM51b7Fu+XqQsD8NYW1d1oSb2cDBH7Mik
uAWxLV0QTj69mkBov3xtQ7F6WUGGg1WzrK79fTKsBnDjbx7BZLzh4E3UGr0o80e9RyDgu9yz3LJD
e33H6e+RRVSmIOoLX+YlRpbTZl50oppDPjm5sHc4hVyH1aIMt/O/UqGcSjdoQc/j1MmSvjpxWsJp
KyIVo5AzWF7hrtb37N19cSBRMRX6xk4UgaasmmGXER01CYIQ3sko4+Cgemi9guMLaC5wcEy4+Qnv
J7JYqb/bau5VlqB9aeQrR9MuFlkrfvPfH6o9XlWvAGRsqBWZ5Fhcs9HbDBKqNfCT0Oq4mcywSYir
cNX9yLeaWCtx6MP+OcRG3h98ct0AhVoHXFOMieliHbGrM5U5O5gTCpsV3+TnPJny5XydxcjBHl7l
zL71pUyBN7IJu/A7myh9Q9g+MUYdAjIDmW1ksXZUjsboYCZ2hWb5dbB54JMfbQHcyQI1e9uOmyTt
EQw50+wELXon7EJdc7NzrXAT26XMPAAblwKwsO32UOsWt7nJGjAKQ6UXpO05vVmFRNoDKgyjw47p
atIrAVmCMCJeZOPlTTGKdLq6jH+Y39YbwoD3I66/T/mRl7Ao2WYTVTQwsHQPN6cNuVao2AeYPrcB
6XveqaAuvwobw6x9t6tNQbdqp0mnQ4tfzPbMCUD/qJU+OTNKfVwuxAJkXz8yd4ZnquLB5p2RWw0R
XQ4APOUVe8kFxPVif5uln6NbkfOqwzBkdhxzPocyDytE/cyN44Z7tMaprxPyvNKX4JPEJRY5J701
UhAlKk9jLzZaxusil4SAGfKaIIpe7HEezOT/6FmUh4Vn37h62eLJrI8M5IfQa+91dmuPOj6PicHV
OqOf2oO2NJa86GvSYQxNHU11HfCP51tn7WJmMJZhxL/2kThjgjRJlcDhJwFXQn4azteSvedESs6Q
KFQt3ZmWP/oAToHSXnkmrGHgGvfkZZSO5JbvWV+rxmIrAGIfePbNONHhZ940k/SY8GTctz+HL+1Z
ytQXP0E3ZPB+NMYz8ZD0DwdPa+Ibl4KfZX0r7W1eDw+a+GQak1ebqX+sjs2enpMKdXBtuqJIq45T
60ub3rWjYS0qoau/iHRbCiqhzTyj8b3Lxw5BrtYdKOEjAMuoAh2S/tjYq2Cd+PfBxPIZ3NTz+8fq
JRqQ/A9xitaw4Hs2mOGiZwJIytP9v2J0ZWUHCsu3wD+0XWI6lRC4wNWCdr3UqdD68GeAVFoE8wls
mf7lbiYUaS0Yp4DuAj+8F0GrsQQVj9one6ChRRZ5K1bzJw6/JzSA0c+suP5i2xNqmd2Hw2JdBXnB
NpuVpOUO15yvq0Yz4BcPJiKGpSzicyMxb1Yw8RJGDPZs62A2KEo6mKbt92cWCuUR8MhvzI1/zIKw
VqlPKhlM43O5rzNIAMOvr2sLOoa2tuSCnb6GusQZN/Pn6Ji5MQFRPpsmrsWDhowa6ZvCMvfu0vun
uA0KSdP4GRIRV88pCyQ1eY66Pbm2xWqF4Dsw1rMCKbx2o7R7gZsI+2mHT3B1RF54/m1+HA3ZU4dt
PvoMAIIg5M6B/dCUKyucCMDpEzY6pGsKCtr5sgA5cSTUuoPeXpgR1vYeWDCrQ0g1oF3ZQ4hJe+v1
YIlL93/vSkLz+4gABHhH8GwzP3TsS4dB1grx4AJn+V4K9OZ+hhDgHaQoYaHLXv9t+mWixnulKlYX
pamklTd1JCMj2iEJ959cKMOgUPcST5GaupIO/Cb0J/2/FAbxQqKiDrWkRW2V1hr06UKFzvOWB9Dw
YhtVNhDgphhdYrTHpjZuFTG637R8l0z9jDqd+lKi4hG+GwlMbgLLrAj2tyYJqJ+FDZAzVs95igfI
9duWVbLFLMyK/hNODFgBtsQMem6N1vU+z/e/Z0nq7mBIAihnNlowG+Nv85RDhOjGtEn6Uw06W9y3
WWiipXflECbULWPEHXPmTSMzgb4PZngF86MqZM1KzkEa5u3GFAyFhQbnLKCgNA5oSXXY682eavKQ
SeJOHGxsg94plAO/mW2OD1AliDy/eh34sGggVyb5sv7qeipUJEwZByAvj/SWlJXlJIF8U5vQLuyr
TMVLGwbdEL611rw9VGERUTl/GR5BjxXO2OmezbtVSgYYE/LhT1U5BxtLGMZjYPdJx6muUs83nMDM
Y7GPo3MZcFX6peA8DEbjFuMAikLhtnTZ8zSH2dmhgfUVV2WJ7HRYtXaxJczmzqdufskF4PYAQOcO
qVSh0fKQo3DIixPNjGBLcE8ybiOY72qnqRlMEy/PBsSSXqPC1kqL/ut+N3osnPyMQTgqWeGQohkK
bwblgt5YwZEdrnynEMzOED/x/e6UEZIKARwugSFYqqjUvPK5/ElY1E4H6kKUj+B+DvAwflqx5hEU
ooWZ7nM/X/jxkqatrVj/1LR7yJPgE0sQwjHmqhr+tizmulZGdeuQATz04lCjt8z9EhhEbcQSLalj
Q9XkMemJrodAQjuHbVXeB4FLi9G8PoJt1Eu7dOaLSLrRZwZWk0KyLPNjJLxxlHtpRpgrBquymxlV
ZgI/Al0QdeUj2RMiWBIHyeX+3lWQQyLeASv3UF2RN9ktshjDVGsZi03HJS4dpV6f/pxcilv06kUE
9fh9tISRflZzcDY+NwcFcHpWan00xFUrC6W7disVMsRDJU/04weeyK9Va42cxHKILLjWbI/QDUag
kJFINXVOMp0iyKtqJMVudr3lInQOTTv7kPB6rUJYniqN3F3S2rAy36ZUviyojePokuvAp4q7NOUe
c1U7m1G4h9gI2g2EuqXdUsMrFJtp0C9q6JxCUEuzgFW049mXtE3HvjU4gBtKkVdkFMadlaJLON/q
Ilms6umBLHvds4oqb/ZgcUZFCHUDSHJAPcEKy8+W+hTbtBHwU+QeOBmRN5bAJKAlSwVCGLCkrS+2
2WKZ4go1aRPNqO2Av79787hm+yguwsPhURDPIaolOuM/RYLHXLOFYm5AubWqHbxbdeoWTmcfEIj5
dmkSdvsktbkYxiaLO2sGQwit38Oqzp/mD/koa5Jdrs8MHOBKREJeALqSB/p08vQFYtzlBNpCWdLp
ltJQfOUcrHXaP4lQ+wAJfzvDSdoOTQa9Q9eXyaVFiKQNBBsfD4yXRAYa6e1Yti/Fapm5FcIXCcWg
D0LIrIfgAgH55Yy3pm+1tShgFEtUjHPsoDMbKyniRCriQJk3eWaz4T//LuM1pR739zJlwYo/ZXnF
TgRrYbva5k1kmThvtYiwgVjHQbaDDrruPpeb68Y302krxTBnFcfNEs199waBOZe1jwQS70/XeDsg
+5yhgDPirttZbKowuXSCymCWXB7p0mz1AjSltDYd+s2FwAsoVbAdTKYAyulKRjglbyodTFUfC67K
IvouEV+dutXcNqvgaiu6I7hKJvgNb70F2lp/J7+i8p3YfL/or+Q3ut9LDmKuyUbM1gcz+UOPJ4nM
Y99twtzxyDEMYTlWfULbDDBuzY6ec2YIN22g/Rdgz6QjGYjos1dbx+UfFxF6whvob2xGPsPlQQay
qDcgsnFimDRJn29ZmSnSF4TNUGboAdt2MAFh2bND8hsdzu3ICW1+mVUwDR89Y4JDMqYiHq0gBPvj
QQMlEQL54f+dAh5RKv1EHyqI9Cmek2h1ANRscaU59dO7sBCaf3cAoFSN7wi5L3a3BF4T+A2tAvfS
/Z7ANAoyqia9xcVJKNnm2AnQS7aYy6fJ3p8qf9juGZniWlUVKQMNgXhFb75It9Gb/S+Y3t0iC62D
7ZcJvPMLQf47FR6E1xg03LKxFbYCfMoTo9O7miQ5tN0RUKVBHMxhNhoQ+sGveBbxqngikOnDIBsW
1ahTs8T3ah6HBAznNug48Q3yAddYFwHWOnGNtbeJ+UsNMIic29u1ILh6jjx0BwUuMVDb3AbslDPn
hGHcNO2fO78xQS+v9Wh5/zgHgh37XlxOHelgN7YBdLYM7dBy0/vwVEqlzv9nY6ju2S97ftfUFVFW
n2NJhizw90NgMJQE0ZT+tKsDaIMmFEBdxyZPUmqVq7drJZMTArFrmJ3IT6QYnVuiqn4XLwnW4V7R
s+xusFXVI29DLUtyI2XDf2GEUIyEuteHxcHYs38AgMmwbkQSHLpM6UB7BBIJL41og15+f3mP3ubh
c2I0ZJb7pVzfmCHT+uevtA5UISPLjOj4csEHN8hNuTt529jw6XOq6LTgBgpTq5pYREOURmlw6MPw
TyKoq/X24IzvLLqRXkDY5cKTWieifrYye1UnmlrPq9PYPMbmLXj/ZS3/bQjWAsFL1th/W4WCGxtJ
ccb4GhvdCT4j3F8xH/x/wI0NTbXGFsYu3vXud9qmD245OTwO10yn2yREOR3UA1hmmK7bF2O+hP4H
CQnqEF6iOYkm2DLs6gTBCv5Pe27pVEJeRF9uzBQz0FSdvUvdq0PRkP0XmxFeykhddGv6VQobs0MU
rY/xbw1Rm080lzcR8OCyhdsx6Sdhq4h3tCqkqMBqaVaLwBhDhXp01zTXdZXoCMfwWLhg7+83DQgR
gRZv539mB82cXGoyEcN3ArRlN6ZuufqVzTHntwsFPKYbIcqi6764zLLGm+2ORwtj8GAiGLqc4CaG
btWQIwcWwgRESbSpjSbakXtLcvgLENF2A7PQpoElCySlQ4ECMk08y8hfMQ+ubm0KZDlka3Gckkd1
HRXKvrxF52R9HLe/wIrnB8NTJiOI95rirO8lf9iplKQyeOCLZzkEFAvbvSc7xzwIEXs0bnoFyXSk
N3u5sw9BtBROhGhKFvbjH4j4Mq8GjL8zpdxeQAB2Wpg65eM8Xtnq8jGy852ySSNLDwbSMUUFnmwY
v6aViSg2tUjAyLJ4uDOuNk+8jG5tAOVGAA3eAU6Xgn1PBwdDqhfRK5a9PRVaaQtYfwLK6sxzRI8i
tSToRo1IuebnhvcaOa7g4tllRd5xkotFcp/8ocQcFq0LuVRGYqYg5XDdaRoYqc+sdOf4RZjrz2rW
45TgueXZX6ukHpHC1GXNc9GW8qG/4a6+rSVK/TwUqJfLzmDhm3E2TjbGmTHr0EZ7SQKFezBAJivO
TSb5ROesknQwYylbgOL9MGhhWmabVAH6p8MQXlk5Oir2hAiXaXgajTKULKcskZMg9+Q85M4SDU4w
Rv6EM6dreA/YHbkdJ9cBuIvt3+qiSrpfgQ0KaVH0ADS8OGHr4XDfhmB8u5GRj7eIqGA8rO4Xvi0X
Zv0AowMA+uS5nwltjp3COpen1DB0Tk8Sszpgh8GZhci5UzRBjPsL50KVmB+dG4BbZJmtOPHLr8xV
8xm4P+n689vUR2H5og5oHH1SX67coAo6EIo9Iyx1rkOcRvPKFMglYBhs6CfeyB+tU0U5+izjkN97
kQfeHLKqLTDkv1ikUVBMH0TlFyUt8S4rsL6KJJceSpgldBLtIvA+1lEprKi6Be/VwIIblT0Jo3MT
QdMQx5Zpg0NEsaaYVOS1OCH01/+tDdhUyhRkzRy040uhhjaLc1dsrnhvWg2DTMF97VzBFPB+nRA9
9rXZ0kOcZNJ8QetdP47N/gPo4UGlLL7Lq4orJiAWLPtPwBxnQ7kVe0gVO/rHwZrjrt1kJt41PW6A
f7s6myvrvmF8/kx6ChDjRkbAH/2Zx6hEhpxuVaNDKjUEUgac3tQ2P7AKwh3tFaTUObYp8SBDEQhI
lA588u4bhAu6YYpezGAvcG+1abw+A4xy9XbTewGSX4xMPGGIq9VIpZpxe/9wGjUUUxbg0mimjPNJ
mpzBcSnS+qmGF5/IhdfOJo+THmVfRc6reJGOTd4qPJnNE6Ogp6wjwa3kT5wPC8JvuENCLm0zgUhz
R2TsF2xrpWIx4eX/aKGWa4wZbULQLR8lF1XK82oK1V0qYXhM/Koj/yv2ujSKuooreH0b06Mz6fdG
zUmasobcqyzM0it/8hhkHBWz7ZNFVt9ecaC8EdjDVAOZHe/hOgz8jssCkhHSl9k/qSBns1Tk2iKi
gEhyg2aRvJg6xTpy/KYK1kmPujrHHPW7LPkc5L2lA0TmQca3X6B72LF4N4P51AUFoftYApF4eypZ
XrhmWYlFCZkBs1A3riivlCw/Le8NVebWBJbi17dajmXym7e8RFN3dLbQ4rwVuJDkUIBU6S3RCuBg
73uFsJtpf/Ts+NJi5MiWMcZRT6JL5JpfhSGJIXi2DdE+pJFjTc7P8lBfh0hF99w3xHcrZ4lJbhfa
PZDwET5yFjpua+0dTjxbSDvzjwtemb3fKB/c7N4nYIvhQ0iM2Pfne7D07evwh1WgNSGppmlW3gvA
UKHgVU/2hr2Ig1s8CHeW7pvsR8bJ+UZlAF+zuT06wGXQy1RaceGiwQd+6j3dnAr5AYg/KWQkTyKG
kdlxOVB0VMxJVny2mFEopRRcSc5TvvDjR8nox5caVTuOH7zSAZBe8WTSLqghLNjC6fMqjbx6cpWc
bzzumYwP1YFn76kEO4JMm1p2yk+2YV8FePQCWuf83wa7KiSRKBqJCaKRfyr82H4AxDcMOm/A1TGA
bhAikDhuTZR5RdKjttTxqISHQ1bvoYmmagS+sTCqZL21PA7hQ/aG9MxuQyq00h9uxJSxGB1x3Q0X
FqWtCO6PmwndUXvV8db2E5cJHq80Lbl4h/C3VKszJqO52BZl3Q4V9zKMMn7e6mFIU2BRbU2mZmv7
z96s7KV5YbCXx+rV0pX7L0qhp4j7HnZoH3jbQhISQw8jHViF6OaX1IfeCfmGSMLae+BoudawweDD
A6qWtLm9CyAAfbyxa6dnM31zMfa5bE3mgPWf4RlTdTbRop3zabvR0+a3ItzmktKa8zZJoaiSL5E1
uWbttPkVc8xhqo1S73Ls2QsMmoZllr7i35f9MF/4h2tfOBHTuA/hn2bx7P5k603EFvIjGRmZvX6m
JvzGsbZtDwSO0Av/yZ8shG4rf+Kffwkl1pkDbJvsBA0Xa4bzDCtRs9wnI0NdrKcRqIdAtgFNs4un
eFWGgdeMVOqAdcVMEcwmvS8etPiULqT5wp1ulIac1dcdo6b+Cs2dQfLQS9R4Ml1OqT027ZrSR/x+
Lse5OJQSL0WN+L6Es8CzKpDDkOJShlwDjgvdQ4uWGxfJNQHut+ihRT86cO97k8Rnq/sh61WXrdfU
4DMI7Z+N33cVadVx9ZN6fTenxBoWLgkFJmDv5fff/EQh1ajtssx3m/iLFapRk3CkboEi/DsDeonC
JURJ3DKTUo5R9wJ2pjU8icc1uWUU37Dv8hTLxkBZwbHOCnXc66ZRL+N6QRgqdPXo0fO5lugd5Cda
VQWyolq/QZVw7cE4C6znqGUOYCCKNlplv4X35qa/d31cDI9D/lfhyG7mInmTaG2QDkA2YvFhe1Lf
nXUFBE7Gv3KwQDv9hbDSG0v9M/7Uv8DBushKaX4lcMNh5KCBu6CSldyJ0UsemhSQoQ5T/x42dyrO
6ZsDaz1DX45d933NTBZqd4qo/zwWV/7pUDCeDb/QIR9g2Lh2PiJwaH/89RF6sh+D86dZfl5JzkFI
9USaUeCUmB4N5+hkZJBU+ukTYVEFL3y3XQ+PrlZ7UnfEAtrUyoN7eKQuX3Szx3Fo/+P2Z9RXnIRr
If/squT+Z/b8vQALeZ2esllWQ6jjWpa19kg/sFBpCOGeT4NGxpzCKTpHKz/dysJ9p649tu35+39H
TxsLCPQ+cNr90DCb1ysDqrDYbCk5K3jqhXJAR/vRMbQjf5Q3UcOKn3G90Q9peM2GAVQ1eEnHvGwQ
yDOfW+7OPNqYRIDA40iHS600VgtCpzFL9ogEsfV3hHgvTvZu9ptlPsIb5tLyqLZxv/Q3q+znQaJz
b+SCdiNsUsYUwRFZ7Mmy47LQ2J+5yBxIlsofXBn3pxOYHJ8A5w5DwuMWMeVoQVWXVD18Yfg/cvN/
akBSGSWjWAZJ+WgAMkMu/eVT6eC7G2woxbaW9TmIdCJuWy8MeqxfHKmDRsmv6ft9qbsisbSmgm7U
ObI5eIHMbMe8quVDnRFbfulVyxlP3xMb/JiWm+KN14PgvOH7DuyoJRB9sNRO3HP4/Po49MaBa8JJ
OHYtiUh91FWi05ouku/n1Tr1o6uX+QYGEyapr2gabX52siTcWiGP17OSE7PgnZ/L7JIHeP4/3QIG
/GuUUZ3WU1Nwn6yv6131jg9YJLFzHgFtJIFWdvr7hDaY59W+BFIWyEL0fNTkyssa2gvnVvVrgvF/
3iuiMEJtC67D2iIWSpBqxklgxGmCWDXkG5zPVWHwp9fgD40tw1ljmSaztjqEN0tpJcovx8hKZPtU
0wulQ7NatSSkN31P7uxKpBnncpbtft2LLmVRUp/cZ/2TxaRWZgCPqP+f5c9paVpjRX7Ylhbfnd90
akat6u8fEbMLTsSzq+j/kAIklbDTqY4A/7U379ypcT62BZ/HJP5qNxxLCOoR64VhZ2Wx+M2FklOw
kO4KSRx34nCNL6g3MQXiC4PqjARnpGWgQi1y7ImU9Sjy5eQA2yLsaCqCgAFn0cXix+YlNB2ivv++
jvry9cKCW+kNmazk24T00a8X1cM5xWgyHMWsgeHPPkQwPWOSXZoAajcE6kK5dGmFLo0SvYshRbIB
GcfJmuRIRZ+rpTbGv0pQ0cBH62wdRJLv/nyT8EChPFRP8qsO9Yf2ZgPxzeHfOHWnjHqN0E0g6bie
hgWkCxjMF0DCDoULWc6FHOCtXHM7ylpEdoeAZ4247voS1C3c+nEYOi/z3C/EOHPU9roqvAYoOaW6
Zb6ll+aiGTMYXGchgQzV8TMIY9pZ2Tlr281CPeOfC6JMMX311akVPEGSuqW4Q8Ya5Y0aCJROYe26
fTEGFdNML7rBdVnKl/qYeWUxkQj9RD+ZxY4C1/tnGem5Y8EB+yQVhwxLOzbdoBWZ0Vh8H4V4uxqi
82K6mbF0u/uRzndmoS/blW19FD5Es5LIPkMmOvFs3iHXtlfZWKZ5BFdr/tvuWlbkJq+ujN/fMOq6
ZHDZNhQCUHJHKUMH+wWsH5MvzubJeg6iAVH/vA9+BrbjKMrID+t+VAzThuAYiAzCIzAbABoA2i6X
TJF7WhkrHoAR6Hu4NYUnH024pejrSVEUlQAD55/Qp166smhv56ublQ/2Da/uEX6m2vsR8aDgVLzh
q49qWsC//b8TzfM0eO2o0cTtSxLBsQeXmm/gqA8d7A0dQqrzT2lVeQKzcfv14aoSnp1dB8DR2xqY
XwQVEO/dnQCErINoTzi4SugAmrIfbeMtAsDbgRk/+YB7GiwfKtEsftkZOJLAWMq3rydLYlH1LdSm
2bhRNah6QOKZ4+E7Uw/RpgvQpe64Fp9/GdA6bKAzTHcuPcaOYHvHQYYFeaXxdM04bQgqIBqSZrWe
qMWCq5R7+jhnCnZLbx86jNrq4GsraCe6QIbBafM6By9Oryx2q9M3YhzxN4dx6vUdQiCVcNtJ81V8
OjOWgUrYIu4hMS+G2yK/NUA+HaNYQv2yjsSOhH/EhtBvrjGiZFapq8I8I9/WY98wa7dgAwE8ohJE
a8xLlce+Dy69w8tSVpmQphDA0DIjEMc6oC1F5KMfPp8QrtpDufb/d0E6G5VtUSJxWzGqPQGnZoS8
1CPdDh3hIJXOLm3lFvQNTFdD5V3ZviNgq196WNg7vKnMGE+6rPHm6R8hRYmUqR1eyV2Q6cunpPQ3
AEXg9DIBoa/VIj9rqbAX9L1lyvY5tvRPWPLXh86twhMf5kJAmss1O9vzJpONSqX0ZNj0Gg8i7B23
dxGbVMzoA7EAYHFJF2SiS9awbVZEg/IROFz6bSqNHz72YUeuR553FJNe+5xtOt57SeanNvlf6+Za
5M/5DaIS122T2CSfPLS4JP4BfjoiPU2OoxTnlrN8O8VNFJ55WqAEJOp6F7kuJCvCTxxQv+hl79Rx
ixcfeWnCOgtT3CRSjl3A0VbVVdOioCs4IeKeBpHLinT5fULn6o2V3lrjThi6LTcFlPmkmbURfgNq
KI/SJBiGZ17himp9Rnw6HAZzVmovDnBaTWp1fljI1Dj3Z/VpFR245H0yda590q+9z/YKfJozQ8Fu
1yB1uW/DU2RC2y8jgMDIgFh9NBbHT0eeR0wHoTiN3LQqifvx6J8yGs7RBgQc85D44p94Y61/YMwW
yRLroKVIhwkNel7gib9sNCHUQoVdXBWpapzRmoIEjDDV3I1vc1aRdrP+l0PiIGhVUr/prvp/Sv+3
iXnPvF8YqDB4J2Qs2dyWzWbMyLAJKD+VL3RUNT+vRH3vHXKjDktU5EFG58/fD7vxdaxNsBZgP9HK
+8msMi3y0LnZv6G5VsjavCKhRipNE7isYpGUYRroh+Z6qKcUFZ90fOmafxCt05pg+I9361uMMnJa
S/j0rYUW9lamQHwd7Oc7czq4+6ii6KfV6duKBfKY4zm/X1Cx8tdE6cVpd4ceVIdq1ubamiXur2mr
sgGgyCIpoSIxuxiHFdE/4Z0GEhKoDuMoRDq2NLjfrUH9zPyI5MYX4suvtAut/B0jsnPlzwJLtmO8
GOgjJzoiX2VTybZXXcDgqQUuiAtPJvK1wrl8kjqlTmMbOWse7lxN702bJAtHBjw3ee62WjVOJx4n
D7KrBWYqTTvuOXez9olMuiffSJTQvxhscWqHmmTsppUQNGOwKn/1hWpakvHq5L3pZvi3fcJtoXzB
VNo2LWnQBW8lcD07Z71+oWo0ytGEzzXE0QQ7aUGdKAEbsf43f2/nZ+4yV/dx59EhcOoUmC5nDuy/
cuQC4FshtkSonGqXTjEVTA0tN+DtuSa/y177mwnmetbKhH6omlq8v3+iGTeo7B74QY9UeG7+xfkr
ztMXUXqt03e8fmWp+8oX2K4Yj4rzX79Utapg9MAfD3F24UgxQXQCTbRkKNeVRshak94omVPvDErl
nMBJ996iQLHgotA1mcXsEHGGrg4oDjxCkfK13We50stfr1wjQbxRvLtqVlH5DDgAgCFWhzsp1IU2
3ZXaPLTFpcunm4nEItc7Of/66yAUcqAH1fmgihuMJYuFbRau92Yi2LO8CkYVv0krQrmtcett0EbY
U5DcM2rJhUZUe5ewCkfcv37TULqsMPgEpUfe2EAuFP0qWPFs5PHl9JJQPqpkvrqf4Rq8zVnpiNZN
k17eHEvu+FDpt38s34N169DTfNvCdjjeTNzJfJvZYbIdiUn+ukPJZCdXzVWWrtTfhVTmNKOz7sNr
fad0NQ1BvRyQXaWGVdgwwFgZos17mBO9zCjac6kgPD2ffxoNElOoWRz9u/Hsktdo/+6U09y8upNg
1WGMMzVFGHMLAnFKadzEXBXrm/I9UeDVMpFNy1NkTSQLpMNhrEctWfzJw6PQkgeJuMbRPDZ3MnsD
9gzRazL0utHKP0j9oMprPzRiHa3xjsVJyr/ELQSAxLao/FtY+MrExPw+1icqSeep1jB9bfC0C9sK
fkY3+YgQiBHiMa0V4ItcpVToKhiHpPiq4GMZrESZu6iZxi80N0yysqXASRJZxfSvvc0amBuY118Y
siNgTJCnvoBJW3nzcUT3GvppTSTknIsgmI0J3t3a/U+2YDl+mtuLs++G9agNxXLc2g8HECjpUoxk
DtQjDDzm7vjItZsFJh1A2jit6JnhSot4cETpF5cCdUipsgl1O/26+CKYoDIMP/J16eXB22QYqbRo
c36IKbCJDzeRQ0z7IUopTeC0emIKIefXqkxCegNWNxa2Gf8t8roPSC9ZXAfjCj4cJHYBh+avuG9u
0Zy0z2E3GNBA+3CXirMvzphUy9rBBFpFnIIxQnXhO2YnMkzo5a5RF67VBeroaaTnKZMKDT/CYUqS
HUrmysoH10vrpzBwjMzv1BiMZnodMCW81+aG8WgmQhOMxKkL4kKQfIoXMmERqIoLtMVKa4b1Qa5R
H/P34i/D17rF5J3s2EDpoCovRm+StYOtsEeniYAsQiXLHjHlJpZlntIYoFdAlmOCYxL7wooiD588
9VXQHQvZA9vNVwuf/+Tppl6MdZtzi130z+XUfcEfVF4mJMT+EJ+vSZ6LBS5ok1ILd0wz8xfCRJzs
bW8oOYwmVGWoDaqmbYA95az+mHQ1dC4CyJjMTXkmuh/GEZMp5cMrctjbYxO9HnvxzblHwLubOv/P
/oN3nTOpL+Ee3R6RxvZHwSvookAsbqhUhyXTrSBM2pnv3MeeN4e/sHQ7fGXjMz632OQuWUYWR8gG
wof20PdP9FJUdfX969KFR2RVOn6y7hC10CQrl3HX9aD3xra6nPd2xW0gzWjsX5dg+DMHRqdGCbBg
X+qxH6U2r6O4mP1hG50HJIScyWdYFAS7BR7xw2+k+iEpFAwhBYxRXWGX6SLysALpgViU3Yfu/8P3
F4+Z6GKG45xj3bx6CkYP81weiQ/hYW3s9jGXsx6m/dirT2ADFskHI/kKeqzRrD8iE/nWM4tMOgGq
iVxNTXmVEforMgDLk8woLmJAEtCWlAG7KNGyqVmVt12vhLQVpONKv4CRrA8mDGNUWf3RsoZuUsHX
LPVESyI3pX3rbHkSKXnT0CgXiObVmVIISoNYo55bZ4m2rSa7CgbRZty658O7CQh+QBBVUUrKrs1r
2NKNreG5mlDV7ca2Z69DujXVqEOcqY9QoV0/X+aA6I+8e2PRtYxPxQR2nHv9vBa5GQUXp3TS50Jo
haUnSGUz7hcBfXplDT/4BDTnz+6Ql1+ntP/FzGPkNsQtlOvnFeF9DZQhva4ZiMznMhrbK84uubc2
XdyG+dK2TRohoZdriH5rEqP7uGLOGMNZZEfuQaGWveXSzYqf5eq0j04VdGyHbCwkbQknijp6/wgs
pn4wkljmDE5FAyK4+umQMCpp0yWMwmGFCcVIDG3d3L2+eqxKSr30Wdbs2ZaMCJqlIuq34p3dIOTd
ljsHzln3ZgMvjZouT5bhEjt6BwY7WDh2zL+FZHP64IrKqnvMHP4TmTtE4d0w4rJIQGyHIDut6b52
R+qXJBkMIrnVeae23RKgCbxagq+6yuqR2NrHKRlB0OputIsGxBaMU72okzuT/Im5c5MY1TzpUTww
u7PcoZSbukNZ89zfsxxoKNizbGuHSR5VoTkG8tt9+dxC4nAUwLWk0buO1rd4ueV0PdT04I81EnNP
xW67DvGBm++IIMQyJ09er0HOt0IJYz1MjRbUgM4HxqukUPSPBzQbElGMBc7rkfZyogRzxArdmIcb
alKuat7TOp2Fh6KkQcskRsl/YZla+n+xB2LfAJIMX8kFhrTdabz8kGIdhfcSwwCppjcm31TDa6Wd
lzssfRZO0WM1pUpH8o56mWqDTc+V9d2BWrHSng5i+Mw7Liwwh4gj/bKaEWliICMQ5l9uuNoeCfiw
kjGYl2CkmoQSHeuFJH+XFukF8a/YeNzHJwMTBKlgmpviDC0iFMRgI8iNIUkPKonSzGuQFDo3PyaU
FYF/DHm5pqkiEMI20VHwS4+/58Zv0d6R5Or8fSXUmmJC59Jzkk/k33GqR6pkEsfiRtacfJQzqw0+
WRdxK48zT8DBoIgaIm4Y+CQaFcUDepBPOSWN+cRBZMdNy2eUrjoLlce8x4RGG8C1BOOU869fF7UT
+vpYUhuS/VebY2Lmsml2h6apU+EmzmbA3ssJAGax6rB5gjSSEr2ws2MJEjHhj02zpCE2NFvAaIcE
PcxJ3PXokGEk107zMl6t39mlb9kYDZHq7fxSA63RE3yJX5zEGQF23JCmu9hpVj11DRncAej0DKCC
DneWUZbEiapRqoTVQdMKK0wC4ovYMsxxo6uJk/IDYRCsgy7Zjq9UGZ1pElLPhWnlEHoO3Kazdv7g
RLn62qQOlttyOPVdkDGIRn/arouzvd4ywuQRIwgb8PoiHTzm4kmTPGTWSgHoXBOk2m1J6O+25e7I
UCaDi6vYqSBsx87v4nRoutGhdCAhTMB+3VhQoT5iZz+QwVQMYWXn3FRJNL5s92wnsFcIrQnPNs9H
5tb+oIZp0Ju6040SkQDPyLFQLiD5hnToiJTz75ZXFNhLLiizlpmkM7YmbYfiPjA47S53wqLAdBLq
kISyQ9EJg3Ke7FT/8bMjJhtTn2JvW8iccYOKiXfGnaVFzplE/mj8e+ESab2MS4lJyrroqD/9wFS/
IyiDbEqq0A7V0F/5IaZ9f/mZroi3PSzUBzvbNuiq3NInApMssunV/qgIHiThFQEbNqRreYiTuIoM
0R66sH30JpZ2o2uqApGty19bKCoVADBderyp0eWrmKx64oiIl2ut5FnpcMhADQk/q7W8Qf+esh33
C6IRKJD5zSv04wnJZJtJxu0wYGCqd3k49AG/BvncvRtuTrzt0DGZFk9HcaTIVkrI5I2/IkfDPues
A4sWRwjGQquQ5KbnVfO7yEWkiWnYJedcDYJzFnRU1/C5Fla2fYYMGZPHqMpAudrNoJ6vCliLj0At
3UKTmF6IFICk5ASmmNpG/T8WBXsNUvsdxAwUhfOg0OIy9ai8xwR7g2PV4Jip1O+W6fz02Uxgqg2r
kH9/kZXLXI60HBAkgzL4Ai9SRQqSXGtbra1iIcoI1ZImob5oePPeSD+HLoLe50jxok0bayPtAkb8
9RXjtOEBwg5Ju2r++K/mVO7hq54R9uTzqUcg685H5aiHKDkVm/fIbKTi/rcVA60cPVxmF/VPBe+e
sFzXD3xHX//AHqteN5lDe0ufjCGUxKDZB8dpqnKahrwjpPx9PZnPomASYK2gzQRPCNbHEjmwbicz
HBTNgQ+aaUy0yyZHcw8DwGyoXyFq9lKMzAHJrT9e3KGqRaNXxusQUkbO5Nhd3bqACNHMWU5gYGei
R5YHPh1ziE1W09ZZIl7pEe6K7lpu3whVQQBsiOXGx06eAP/r8BBHTOpLrsjW2fNt4pSI9DnAzGMY
4eKUnT4WL2Nc6ioeUFlchi31PyJcd9Qg82urYrTbpLWsk9bZxqJ4JC1dNL4GQ6ZEe31umpyHV0jq
Vh1Pb4Gti5jY8DCLlQtAbOHYZLqcIk1NBMjkxs9QS7kJxI8vfCyMreu7GJAQuI+tEZaJkYu8reFi
A4abJ5JF21TKUnzecY4MxjFcO1l/8JfRmeQ21YiXgB9n0fJu+aETCOeMjcn6wnOzU89+EW1Mck9Q
dZ1c3lli1b2ssdA4IgSJ759N+ZOguGjW63GxdsIFi4vvRgBLmtXtcV1+3xqoZwhLDnW71qFQv+YX
/Gl9NFz5g8PnzYgRJ91vIzC0tWxYxpGhW178pXOouIVH6pjeEa7ws9VEAFPyHibNFwQ6d+O75tcn
QHAn018dd5XXCx3IcW8L42IagmsTc/6u4wOBAtIEMMYcKnesTiXoBaMapa0zF3KT6oh7qeFE7FC5
uX38rUggiZLAfU3s/t4mh0vtwN9Xs4Mdh/FcBMexcsd3z1xAAUzueKeACeyOYvkFKMA6vCqBUI6c
gnAS1vu8WO8uuMwEJZlttT/UV7Gg5VXtPPtKJO3ysFOb9EfTQLfbFOSYecVNnCsnv+C7fstebu7i
XMwIFpg/F38T1OrUChcKbm4xCUeczMa7B0Wa8c0k7Yf0bMDRcTF4ywhK5XUGXi/O5wr+i3EprvkX
+oH8slSnt4BEsvoFa+zvv1j+NVAM/SEbZ3ukOMpH5Pk95kWROiJ8p+HaZc8hOT+2KLfFt2sTNO+A
Z1UR5RZQYCdXSvYYvCwhyJkwju/6tk/5sdKRw5igZuCqA2DuApa1ZeBUG20ZdkLe6pVszAzq6ml4
5BRddVfLqbARA82p3U0jXIFCAeW0KWf3SZRKB9KCqp5Ygz9Gh4/45decnfTDSacY4/UZ20qLdFNX
k52G+FpTNhosGsmPc6LDB4VkMBcZVvbbQ+JvTzaAlalYfRk24v70X34Hjbp71F0sRjpwMjqgbsuv
eJjD8JWHS6F+IxN149OzoFfbsYTL2o12FQaquMcAx6S+0IuNIkU7L22V+7hiN1SWjGDilHuy95PO
wX7SEdauYBvLFwQIhGe9ubjXyZLZCvPT3UO7SKSkXlPLpzIIEwVX3qzBEjXHXO/jqBDt6gPIBL3U
QhUauRIjPzIhpXi7BrFpxDC/a1cafcxS4RMxgAZZDmfvoljYoabV2L6EnU0jM/OC3qbPK8xQPlYg
bNlRanrTIhzTESmwW1Zutud7Qx1z8UnriCyFWMQQSyZ2VJBanjcBkfm+BOKybRw2BRX9+KWEtZWS
4pojRScCA24CxKZTUxLU6XCtPd/WnG+I+7+loLlsVlQA6KuAln8NAoPxGHUlj/jVK6V0+Bq9Khdb
n1WSvYoIXCI3eEr4ht7q0u3aHbNq0x8dMi2imMAB3IYRVIzov/Xo0gZbl7q40clW0UVQwoKparzN
SclfFnzcsZjvOwsxmrBF/aXJP0Y56JzwMrPkpLq/PNSwttzKjBF1nzXUMCT/Vmmq2ux0/EoxEFi8
vN3lcUbmppqzudY4nXMg+6FATZJ/TyI2PlVungrp3fGVRrSEh1wlAnwl+RcuhwMa9T91HS1P6aBn
slyD2mogyJjWjHxJMbbl76ttxQjGgzHJMAoOBCsGijx/q6unB6MlQbv6w8uP8c4wjBCWs5zc5hPJ
1WYlGxFeWbiwQVOP0BUgeNAz2eeNx9rGLx7uDdXv1eczBjNbOccPtuzQlTvIJkm3D5H/nxSVP0Qe
G52GuacL2qahmebgQBpmsa3PVws75OKBDu7zGZSoxkZue0Tw7bef4ktjcbsjvyK6ghSl2Jo6fkj/
99+1FoMn89C2vLx4fpkwKZiV/5wQmlqW4CEMaYROWWeP9XshLW/NGwYuS+6a7SXDjk+rbnart9ym
0waXri7PqIvObzf05nZSPhkjBJZpfunDMUGRk9BNxEwps8OjygAYaU9ZhZjdw8haAv3JdQ8d+dYY
tjiKQEtUUgBRh2WjhAhYSiOMAqJklan4TcjQzHgbNTgq70HXCw7hbz0w87tyD531BepjrEgF7WDq
i87KL1mWe04o6U8Gr2zp7svLclK7SW/befYM9i3aQ47esZgOZhIP/6XYOhkw7sOVQsDghxwUVR7i
EFOI7jjfnyh78VuCT9CH0Yhf+4bHZ4K01wvEw7kKf1naZ+ZkMSnQbG0QSD6KX9PO0LB6Qz9ZXfln
VCVSBrSLnDHpUkPQd0I9bPJLZhrnHwgKkkib0B5w1vdEdKR8UU0X7cCa/XaMlM2q/t9H2AmCOTug
jWzFGucIt7C1cOU5br6I6v8NRqSI8O02UCVaXGuPMHuKpQe3jEHlLzGk05MzlrPBE8PqQe7PQWcf
uCK4xkLLQexcr27CX9niov0qrhChB+UxxhFrp7BZJyMAu/jigSjANYpWgzBqGIIwEs8w5aAwKinb
SwEmbYLJc9yqY7ZLDUv9gWtKcn9oFXHhkb5OX9o8yCoxeYWXNcVY/0Y1hpxhKXl/OrDysOb/RdIQ
GJLn/WwFPye5SgJz+w9ODYG48fFi7FYknVG9pFsQcXwyKe+Dl+FCpR3kg27PLIcnRjmlF6AWwXbM
Dm97oaGxN5EgQy9SHZ22X34TO1Exxw/2ENZUTlNvxDGapX14SIUeXXQEvnHYRKL9dx6O/XrHzVvN
TQb1933t8fnl9OrSPIlog81af/QbPoDrnOMmLldHv3zwnsCSsn2SEQ+PHN+O5aVypojdS8ZSNZep
04Uel9a6Aw3cy368B/RTS0zfsBAnkQREe8oLMQ+POyAf30gUhNu/NL67ggvC/xHw6+yZ+QPGP4QU
F4swP875aCr+Ke0/pNQKXK6KeH0TZ9wDvdaEuCvlCdvjs5c/LxrVTmQtUwUvkrcAF4w0GzjvzpWV
vpghDFbuwdJNgneocQOPF5YIzyoV9vAuWoDWu+9BcThlX5qew9uwe6BhyzJj+msRyScEmxlRYV12
NhU3RveImhMO7h/kzeP7FarDev83pLiWb7rCXcUvlq7YYzPeRsB+P2RVxuZ2DYvlncWMbz2u0EPX
bwFRHfDOxmyESsLAnrpIxmKqG2cCo/mpFf8jET7B8zPWE31KElINluMRc8xQXe+tXB0Y50pbSK1I
mQRGEIz/i0yhPbH4cateiqbal2J4PR+K10Hp5mqJZwsaf2HpoX2hRvBP5D8F5uOOBPq3x1laVR9Z
nHyWv2KawvyNl65klEOFE2Ub9IjQw+OEB/1tOM62ZE+ZGeVxxtARDhhOla4lDRqfwvIFhVT39Hvs
VVGL6ki47vzxHVMPGPLz4unkiu09AXB5EXUUUwol16m0HhoKkqP1EgjQZxg9o9X6FSUVkxQU6r6c
ZNntVxk7z7yeLg3rJt5HUWXba4FPp/hLOQvz5XFcLreunBhQcs3ooZzG2TKNOrrCJ6u1FhQKec3J
k/u8xO3qExWi69BXXLrbPuMO0Sq/CnVkJU4Zh2ez9SKhQ+hO0aL+3wcWyQsZPVA2cRi+i6K6rl+z
L/XfaKckS0tco+2nPSj935PNaPPPx2ceMB5VvdZdO9oOwTgigBIMLv529TlQD0zz2xSCJISbaD+8
JUItU8xOVHD8Iwcw4BdsLIKjQhdirNQBJN+E4lDWnEdG7ZMZcp6UMidmOe+e7HWpvxSt6SYUIUdP
h1sO3I9VHQmwnLoCCcWNvRClll3eO8Iao/mGptxzXZ3nhzyBeJvRTMWe5JnHwBi/9z1rNWeuY0nf
efVVTugKEd1XWMhzbMuNToqllM5XQ7kl+TXyX2YcthQd1og0HFl6gLr1mwFb3gdHecqxhou0Th0f
Eu2FKuN2Fyil/+a6Oy1rgqR5ZPFkN1Ru1pd001A4RHDN/NViQqr3aF6jJOeq8egeLOf4nXB5W+er
j0fkpvHF1erkzseZdDyKP7fE1LWF7dBkpLGQU+Vm7ljrepGm1WkMp+PGzYXDvCngzWFlkbCFo9aO
uDX/N/8pF8jPeQMHzpcmGu339Cc/5NsyUm4STLgu2kIvvJWub5qaE+iQUtQfEAV2r7QdOTImbCzX
vdHPnD82gIlSncoQAlPoHs2w0vqIQhCoIy53QATHli9CtAb1YCSMcEOaoM0WL7qvfSYwjgJypLWW
Sv7kg25C9XqEvPFow4r7D3rBslGmUw9916Mq/0wpuv1EKE10uwXPy7FUd0lmKjm1VIpuMxXsu0N1
Y4t7YgQDIRnDqPkdxnaHID0mFh2+x+x9nGUC0er5tbndeh/p8AclJo94ICiRK6f1y2Im9yAZVtJ2
EzoDV1izmBKozrebbO4LJo+0MVL3ftmA0IFvaeBmqfZq9+rZWJP2nNXwFvkeM8Le50lZSz4+LLyn
6F4IAUvTCRrBzCmAfISyMR5pd8xRBdqFnhadsQNg5mBzyMRRxAMl6jwg/ugOWLIKoPGZD5kX7KPC
NQHxRvpf/Da7+mQHwCWPQnOY0z5cBcDgeJ/mtsC6G9xmeF2nb20Z0vwQz2ZFzLaNJOJr2ndg+N5S
4ezln5uRL/Dw0U+gqqVJbwmxzV1YIVy8UL3g9CvyC4ilJqxdGeSs/pkWiMi0AyftPAj19zKvaPNt
FV8jmbshUkMyaHCzp5KUg9iCwErTb/JBS8ZcUFw25y2n13v/glml+ygu1yr0VwCfBmaCzIyNtVpv
rMxt2LI9qsVQWhnkWx2q5EqTa92RmXXhW6ynB3LfsvSMpMfsC8kRMhVOT17RHkfhdy+n1ckKXu0g
RL7pgv6w7r6rQCxyKOZ2J5s/VYpo1CaBcT74ytFlfw8dCnKa2282Cb7bOl7xGfGgYIdofCFrqk/z
4veWrZS3Cf83WxFod1UooH4a9PIrkFwAr+M6mPD8u9Iqf3WJi9dtnCD7/0WHXQ078CNlk03a/P6x
YPVXSttcuXFmqw75zXNayYoMVif681+h3Wp0/Bgl5fiTd1d7qcIaggkeaYhgn+rsa84e0Q0bPU6Y
UGsO+Vd3m+X6ZXnuqWmzdOHzvSB5XEL/ZWeoIQX6aRM4GgBMYQZFOryfzDU3zW987jnVGcopb7kY
JXpJtzqF2NQQzheukaAXUrOzbVh1P2MfKQFJFENpMs7aKAXEj88hxT8glUWrVB8FJDr0rWhbRrjw
wqs8ypk+SGc3j0owpaF2BsRntECu2D3EYcdN1eJ9jd42eZJEsJGFi8q+zdgfizbzo3nbcUJDmnKK
rz0LNCXWrk5ZlqylMoTsba+fUOhgdCJ4agtDFLbZxRHCyNc/hSNA5dSbirL8T7Qzx35Mym/vT++K
YrQbp/bRlZjM/tEVcRmQSAEExxoOfJywAFIynwVKPWFApkzsVbkyg0n2BiREfJ5FQqon7l8OE1SL
+mp4YqKDDwie8hyBM1RJyE9EFkzTgEtGCvL7IWSoUjtMZGdYcx/m6hyffv1A+VvnivKPpeHqwNP4
sJSYkq7vj7j7tpIQ21XoziDtbuCRuNn+XLVxyKaOMqZ3JO2VHYjDY5s0wsRsXjJkjnbzYS5R1KrQ
O5XxCIX7kHWnsgHB2X9V7ObK0c8jsx95pXr9Hx/o21a6JeEEGqU82ood7dmcCFDlj0kC0vSOZSWw
//m/J1jga8kxq/onFnyf0G/0DFJk2/AsniG/lWs7nTkEeAB/nK6ErN11uDr2gOc6xifn5wJuCJBL
UCVIav6KEQUvqg6ZVJHjqxtsgeQ1smm+oCXUq9jD/XgCuJuTbn9VnyaAI/SGeve6wFOapXLwdXFD
l9HctPAI+ubQep30OhMT93JdoZZCMmV60oLr5I+QKpzKlQ0/s8IM8eLHxUS5RDR+VyBev9mguz+z
JHYcEd6vhu1DiL1sFOdAjOc/SgjPzSlqXohpglxvZQ43uvVL9yjV0oeGN3mce+o40j//mkWreGcA
iE/S8YPIVNjuk3I6WFwMvgxBjonX1wgOe4kICIIol9tvbJjg+DKqeOcJLPQtbgWzxKHA/HJwtbXd
uJNJ8eiBK265rhEjcYas/709yYg4ZSYkPasnXNzylGP4t3ldNiRa9gtze5wd8oTVD9YKiDweS/uS
LrenPY7TMjzSf7H4oHgH1LioQDY0Iz4gJ2mhO8BIOvNvbNxpug3xWy52ZVyZFrI4JQdTPcWzkGTQ
btjMCRjP5X+AXAGlQiLG0KQnJi0teAQfl/v3HM2YKrl0CPi+ZRJGnPwxv9K9lLJpuEcxH47IUB2F
Oo9z8pNLUEQftBmV34H8q7TiSeR3j2KpoQ8JOwvSMAQXS15Q10XMFd+PnneBzmqkAD64OJic4xEn
1t2lTBjTkGuZOA8Mi3Hnx9WKMaxNZ/osdMrXY9XneADZYE3Ct3Cse2n0003X4AQxCfPlPQg/0LcG
JrNWPO6GYlatO9LM53HYfGQTgn6TALgQCke8MGPXyq9FDJZ5/Ed0WEf923CVLORcjWttshUAnosW
Rpt0Oh1mbNeuvNFeQijyvoiDbDWGDSTXwK5IBfVMaZQyMqMvcq41xaVkPxwnTyVLbb+iFkqKsB+t
FjGUKFplXWNA1KnK9xMg3jy0UampOhYdggWyMZ4f4nmkG6tIpJvVfoGVXfH46OgLyshVQHJcQ2k/
mUcurGbfo7OramAOOwK8MrbFyGObEMGLE1JKmUSYnvueFtEaygBDhSnhEdgtFgDqbgbuwpCKsejL
w1epEqTmr2ClCPIHF+33ZVcf4B8Cj5nvL8md27A1RbbXrdqgRxs0Z9r0Pn9LoL+W2V655F+ejJVf
9noD/J5GxooerZ1cnWTQXQKD7jXm8vP8YkpwUMGs17Lw7m0xzcVMl9DcC1Hucwf9U66rUUhUPfEi
xlgoVCgGecYZ3jtt/A4WTWlMvXOePCk69pDxThiqZLx2Zh5FR3U1QFXkipuHZSeR/rOzD5/jQUwS
jU/s3kXtGHhT+Uvh4LlC3YfTqt7W3ZvXUER+hN+xBnxwpUb9CZHWKaMiwfc13eNcX2wnu4CTOepw
rEvm1wd6HfIhQpO9LCU+3qP/3IMRroqJ9LMVZT4Js/YGJI27eqowGs1dX/njC75Z9yQ3J5NRHm+B
m3WAmjeYGk3aW7XHOT3GNsKR73I7x+TluimhGLX8M0VFaJp8pM9E0YooChqlHdJ+WXVtpUNIGq/X
gJbtdUT53umS6S0fm4yGWtDuhvmswpgWmAeUpTWKduiw5wnsV9ZIoGQ2GeHtODoarOh19kPol/PZ
8XSiO2OL/9hu/OZl7k0pkkTHHsGyGJPm6jgR1vPw172g6t5oQ8NE22Fu9hlbPb//oKLNW33xRFBj
H4mJXyvpuaAHx9U8kFhLCefMTrAr/72m1w+hsFj+gdCh5nbVlGSbxUNGoBDzFmQH3kzs3W4ThAiG
YVfAoxNztesisTl4YrJ4AXmGuaXQ+LhQxwpahmdWu/yjr39vOnYe6VIOAr/WpH83crLM8aliYdCe
qTQsl359qZeUNhsalC2noGoL3Ls9LghwKZd9lmI5UVDVmnw7JfsuklAbYGHuWFOzhWx6mm/XmOC7
Ca4EOO9m74vpY8ceEcOPF0pXLQUEMHd7sbUFBPKGLqVi4NiS+I3aDOrH4ivnQnmV5lQ0XbjdLLL4
x0omUWtPs2Xiis9GUbYLk5S814hJsvf1J30+nnctCUyzMrL/CyfMCPsfx+2TDh7ISZ8EsvgDAW+s
fV9vUd8pKbRqYFkhUi2n1hhlmlQBxaXOzgocFG4Exu4pQN2LbUkstYSwxsXCfzMBmxu5LW11IQ48
r/XSKCuWzLCMgWyTN8ONuqQLnceanz+k2vDdof+2LM0uQ1XbUqmaaJY816mXNIoPwM0a+YhSvSYD
EelZBn5Kc8VpTAnxtrUUOxHf/7wfxSC6UUlDRpumPRT5dIdsly4WxeOnbRh7g3l+XFsPy/nvaQa9
rzUUaC0WvN0XrpBRboG/JJOI5g3J7VGaN+vbKOHGHZ+K+xqEQXKVN7wSwBF/dsul+IiNjYUdzkCw
xKNhonVFEww+jqZwElY5DeArOJNl1Hpg++zVRVRRsvianpmFDWSjUW79eREr63j+m3jo3Rzr2+1b
1CLq0bc+PYhQzH+nJWViQYBKDPMhX6S+vq9ZTugM1H+CiV7C/1jvteotRP/VVJ88SqlwNq7ObbWL
ETLrJZg2EwwlS0rFb2sIDvv+1HBOeSkYASG/fKnFM4fsTSFODB0Ad7uLG5SwL8LtGa1jFXYd7bSp
Z9yGyGVX0oBCCkgKbIKR0zzhOMMJBut00mMVsIHJBquuA+1IQWiGVKjfmSLnRC7Gixx28b6YNLKe
T4lr4LnMN5X5hhMlg2AQzL2QyST/hAcef75TMdomo5u0qXFo33fEn7r4/xMLotps9ZefM5uePYS5
5c6daQxdpvYM84ymea+F5IIRBmU8eO9/53YVgLcx5UxoWcSc7Q3nUb2IAnMAA2MHpRNDOPiul3KB
4cyYA6U05BLqGw6M0okyteqJiyDzzjVk7lN7aEF9gC/P6c7d1dIYqqrDj1CQk51SpVCf/Uiy25Uo
EfAioTUeBD40nJjieZS1bwdF9xtfAx+U58tJF97cPWamDXrq/H2bcbSSioU1B2Tnn/BJB6KI2D9I
nzU/BIYGnYm157nHVvUvA+zZGAsib+V35r0tNKJnjeleJxsMZAn2AaUOSSVpmvXha26asvEpUvo9
mdIKys1WMIO9YcQdx3AtqS3DEFXgOtT01ggDozec1LdmmZ8PNyGVhTnt9PpfxUftO1o/vY1NihUw
KseBnUKG+u48O5btAH9waL61zzYObjaVRCCbXAJLZTHFO3lS4wVWQOPegLQTFSK6HeGQdXlEtqyU
27I95fy/iSbav4ami/PorhscLxD57abxBXBB6E6YYNysipQpCPmt9xlqXRvWX3/AExuPF/eP4Ddf
dIu/FA7sYVmBiaMKbYo9qhkHXUDm87Zq9RkClLqXpO7qyda5ldXd+G29PmW+US3VISDGOALZXPsq
IjDSo1n7MD6VhlYg/WraJ77VJ1DR+gNP3bpUu9GFz206oijsQIKj8G518vjxWC+JOuaFMVF2Xe7d
yGtq2PDUCYp9HMG4VOiT7lALias6Uf7qkEi/n0nxkI3L5230jy7r+8V9TuQJK22gw/ruPnRI/7oK
+QYTBv+GTovvbmSkGLiHcpsNNGwlW1LcYnzRzOyODSU2Nq2lON/AJkqwKiapLKveRlgn1L0Aqp4n
YWk08y3MSDOukJptlp3xkVV6KR48rgABn5RsX2PZt3devTu6gcmQLpZ5TUAJ2cxOfDT6o9aCRGac
mlcPbx+SjtBzy6XWck3Yi4/+kN3yhepa13Z2R0jMTlmHJfhE2OYJNb61EMBi94vqcHF+AY4lgdgP
DPob1StTUGGKT3kj8IiI2zZQScUDbsSbntY7dOvrFLia4Caj6rXSs1M028qYIRbAxgGMKdi5TcGd
RMcpi90v1UxH3GGpQCE8e6PojQe9dxLgg7XvG4/z+eQWJ4rZieoa2ZWg42xawtSvtC/DrmM8M0Md
/jN5eXCMHBZ5jSg8ouJ/0E/nPhyOtfkYQtwxcDbjjrf1o3TO++hFq0SRKA5/xEp7kB3nK7KigwL7
hcgnVPWBAP0w9Yi4IH6Y595Og7hwBBskm0fzGBTlaiZrPKh3eDQs38H337xV4GchXhmiIR2DgFXN
zy/v0plId7JXWjtpI4Xs+avt0U1aIkEV3c4DMyN5E4LEYpmUisjeVk7Tw+AQjhd9n2/B3ortMqS+
msDnGx062TqUl/c9e4d5fMjczBBq+ud2/k+QdN6kF7Blip3sitX/d4tH7K0biAgvsBSEPsNc5yOq
+1bhMNuqnhS81ex4gMGDvgP73T0aXt0tIa5OGpYc43vZZyCvcisUWrcDq3qjcdFyuLG9xGi6e1hD
P9xe4ZapxjQ0BgscRK5N7XNw0kK7Hf2O3+z4ARUx7CqOYpWuk8nZOl4I6fhhDZhKOuUVp/s2324u
G+6Y5wM+20n/qNinIH0+KUkIVfjkPI+h2sXF2AjrnnWxoV/M2OOI4UCR2Jug5+06lOdBVpqUZEdg
6bHMAZViyTzqwSdew9BMK7eacey1yWN9z6NErCkSTwMU/+JtF7qYblBs/xHkfYgMgZJpPxBoUQe/
RY6jt9s7PxVT6XzpWmKBwpLPZaCaL0kJdA6qgH1FZkWmkd56mxoiWbcQ5RBPs59uY4fOCnyE4NVs
EMMOuLD7z7whvDiT2SyxeaAEdkFEowHxMyTHNJobRQEje5EnFTt4VeSKAs8eF+qoORW5cZTeu3PR
H7cezje7txqRqtqK728KduJC7BZklq0tVdf5kBSSPYO0ccc1kQVGe5kur3K43Tzyjn4Y9856PZ7P
nDL7u7Bej0qKsrz75enfaCDqbzfEBpwZmjC2BsEgG+hIHz+KGS5wiwxCyI2qXiqp7/qklbbEz8vH
vxgLUff16c2oYhSKCshE01KcsYTfaY9L7cGCQCN/yh9JZqiidSNFSrWlDV73Q/G2C7wISXLBMvw8
DOKxLjhEVPvuw6WY0DvirWiVdgtUffwuY7+QTY3YxOjIHko9cLi/0m/rjUhqcUH7G4tR2inbkuUe
a5hZvziShc/hL+rmlWRBM9yqpUO3vt7DVQmDNrIeFstV38J5HjyL7BQglhBVMxxLEfh/zrUV2OXt
/qKlTnt9dRHEkpkF4Afvf2GPmub4wBDKBApmTEXUq0y/7mZboMuyl1Kv3DSpcGjsexrrnRUJATk/
RZHtAsgI9cqmdNqXzVbBRkN4gIlOUb1zHtNyjOolPDyy2qaXP45eYM18fC+f3XX38KMPRAqQ5upC
mrl5Az2Kiohw/Xdyu4nbvkbGJJtOljnDoB+WfwKzfik9+s84498qWKBIb9rLMgdwJqH0pA6ZItUo
DBq+CsV7OS4Fn54sl4RRQddQG4s54srkYyF4AT9er58xMNkI8zOsYXCRxAcA3CmrhEtIP03ik1N0
ilau/DjILxU9u4UYkCqrBf+FH2a+NVYllVq9vuD7HFkNgkK/Rmil/l1uBFNJp80yV6fgI+bUN8AY
qeR8y1YksgCEg7VnHPphtQKm2Pjhk/RzAaWk4qGwoGVzpjFuK8hYLvlxeyl6yQh+ZEoK9dymq+qQ
HGS7fL1Hyf0PgyKFN9rY9XeLVI9cLkZvR/1WoKjPHQOU9oKf+uU5kEAZCfIijb28+4Km4icdXo49
tqmzXEnjpI1ABAGTrcGZNiMAIrgV85uLykXp35waB8GaUbXplzkS9su3PR+SV1+zzsWpffCaz0f4
bDHi5rAB69/vf8yQYs1Oqfmd2q9Km1UTbxdXShWC87OWeXnelwgwk2hnWuRHknbtH6CdG6VXJaz+
tO5+FgYNQD8FT4nELhHqZC37z5DS5Q6CZfhxb94mplxxDRgKHJjrHwiRgJHyGW5CVcmEOcRmjgQH
XAdEYdi+pWS/fn69ARQWILbSiHstwnux/0Q8SwYY1M3wzQRM/OQ4+5pS3AHljLxxKb775iCRlrlA
9fFHZCa1986PTgjndMfd9PBn1zZkkg1w+lIZKC3asf2HDIV5TUNRdyV8/cI/IdR+/QXYWAr2wPiB
dXAWmfpIJ3f77bixWFdisoSwnDFpIj3uvF27X9RyvfBQToSVkhIWCC96fjsUNqA9RlfCiBU5rVnR
6Gwe5Va+p00ieoV54XoeuD5YbcoMC45VfOKWALml+4SvtjaUT1W+ex4eUkkcRPTZKGUoQmei6ELx
uNdtD93RCfxizZuR9f4SCfZmiNiZV1PwrlRju4sMaFuo+4+cg8/4U4sPUvLKRpQrwTT3cW/y8YPm
8SmpTZaF+qocjQxnBkROe4X876L2IA7++FJKROy6b+kSscIoGBCd5AsHKqjBgTiWTXuPFFyDv4C3
wyzOQuEIJx3+95GAcDPYpBzCBPJ647o+uPXv2LAsHsfph9pI3cudSwx96rIMOHruhav/beJ86i9J
QyZheypXpDLTEdJ05+b0iCD0V3PvXC8TB1DFSMvMljUfwaZj5+qGaVEFKcT1SZDOlBZNHf0IWWQG
lkif6VcnaJ58R/fI3uH03kpw6wvwC7bLus4t7rlR02fYRXIM+e+c90EhCaPHWKQ5hf8qzHM8Ui8+
Y6w8MvHuVq88SjsA5xchlMkm5mOKSF09kwO3NGnkGgD8DM9OHybG+Hsp+Q3n//nuAnD/Sw109NEw
LUHXw3RAWjsTEExVYRu+dlQdfXXFsIx5V8Dk1hAPVzMKfttUznfiQxHGb0Yce/fGq9IKa5qZPvaN
H1G+M+dJLBcxe9c1DFEpZHjTUiv5qelvABcYUGxJdwLee9H1IIV/vpBhPzC+sgkjxA5dvAOy8NJ5
yRY97mGLxtWmJEoGTHMn9w3o4tIQCO2UcGC8z/a/YEJjOUL0/sOFYGZdnipEAF6P3wHoJkDGppO4
NBon3IXcs/Yrd2M0AGTjeyMwuvz7T/6VzFX9LWFKgtJpq7cukXPMIG30oCtd3LrPSsZXkUiune5d
Ui0HoUxnmDjoymO1+zLq28HuhqooJk028++RRDyCgPLzkiUygIfobbGUhGeCvoX1A6KjPFwP2+Oi
pxvexNuiUOiZRpEIP4FztaBGy2DvPY56ed0YWV8PHKCXtBVJFzErN4Oman4LFRcCup21WpEtbUuQ
3Cc8Xx9H+QPwth5QWHD0+NGXn3K4tqYZPro3HWLRKf4K638gF8LOotQh6t8YM3U521Blt29MVD7g
owPPUsTkvMgpL5iY85GqHpRbMAldPMhG6IGtWWGrxPM8RT7NeJt8s8JUQiethRuqgY3pqmG4/J6C
NHjmmnEn218/iAkT32OF2CJAMV06GDp8UqJZ55S54GkUVZ+7OLZUNRpK+QfXJQdcErhmqIJCzLDa
lToNIUCR/2JHppxs2XBKp+zwmv9xATAtqS0vJ0u27N3bWnM36mxKbh3w6gaTknuPqDw3OqjW7oE5
4pIM/qdj1vlk7RmDurHb7G3CEQ4/1ewQ/cz8DsUw32zcWEQzJ0zfidqwVZgx08lIoH8gV5Xul+I4
Xb6XR7bNgB5LJIC6s4ANkzfJAS2MOuCftdLr+vImuLA+Ew9fBuCgQIezUU/PMPdfCixBvljkSGZm
w5mEzp+NuroLKJc+HIEZ4GIpETpvZ75H0Wr+hvSKn3QeLuYGJjc13MjzghMY5rK/oj3QXv2M6S05
tsymU7mCO4IcgUCIW6SFeSH5Y/hAXbtrHBH66LrEvO9rujSySl2nhEPDUoG4k4V3voUfdesMTAY6
ORbIPemj2FeoeT4/vapAh5Mn9OXLTEXhApZeCVerw07BrSOu8NhZvlaHdWgv3aYZfYfurwd724TG
RiDPxY+rF9iX8dpsC+x2rHypyt1YwCrq33/ReRUb4IQe/BEGcBEo8FS6hkiBYQJEIx4KW/H3z3W2
EM6L5+FSW6PeHSbfid+Qdixdt91AREKt6STTusUgY7M0N4C2VFyrwHMzwVQ+GOrpOvq8HMtGdEcJ
phLw/myROZ+u7jhqn7LkSzTjZzvqYFefHLJTMPFfO2ZwKaIcbtXCk6YnDwiPQcKYCCzhbgvLRjYK
g0JI9/pUVRxsGlchXcLSpaByRJMsC9knCPcbxp+4fuBF2qaUA+c5EO6rRa0s/zrM8bhqaNyDWhbH
w8F6+viXHqAW6q/+owQSZMMei0Zl9zVT19g6CHjoIBZe3rZ4rCB2Zrz09adC3vVjMcWx8wkjVtge
q9YQWXK9XWr5ZeT9/BJ6+PHQMcPKMDhWA/vhtYs/mnFrtIznFz90tgBuB79DbYL8Vg7syW0xE3Gw
JkaWwxE8rZG45nQZzSaoMYM54WkdcWqyv0Apzic4EzWgk2XuAHczizF5JdhtIhAL1MNZm1gyebo9
7JgC5pozksR2wo6dWmHGBLd2Km6zlx6ebVr6GpOSs4aLH8qTXn8OqxT3jkj5ii6xW5RaPv6UoMnV
qzDiPVU0Ohm422WVu/egJPRoSWUDg32UdH6R9QNLpTI+YneYI8hYbXeH3rNLzu6sTzdCfFKk2px1
EOF04/FWE2RlOitjH+RLDiDxXtkHLAnpzaM0vG8px2GNg3B8U8rDbsjVAztgRdxjFnz8pVxO2Ub8
TBvyGdDcXwAnbX/Wh9+X+3uB76Bj5OZzNhYWMHWBNwDh8dkK3zXgwT+WOTLRW/PAWyR/EMakHBtB
rwBsJzEcXI3U0MwwLEsv+Qhg91gpYY10jTsbkymGyKCnIHDuU5MJfESq2e7xk+hmKnvRzsMTCUTh
HtIo4hAVbko9jdAIlAKSlMeqOIa21wqtI83SRrXVUs1/OHrsr63CLrK3lF+q08QYKOFARNzkRbAa
jHM5xuGtR/4ZIJOp0wWDa9C7hEIyqJ28f1ze84zb2fAJLGFD7tT9MjPs7Fqm2F9Ba3LNVK6S3BBw
e16r46gUa+h0pB2QkTsWEhGJOvayfWqsbL/s6TCdy0v+QN8p2wUExBlFrGyO0SZmtu9egWiJzPOj
O+xqwhcdXtJofa3jowiwhq813Ae5Dc2/0SADI3GtxRmo6xPKHLkHBf8+9ok7Z385TnBKMmhDtfnn
M3rMZ0DlNhcjwD/yqcRQrl/uBDDWxisgEOHwUc7O2QJFAmwSwb/Mdt6D8UV7cfFGFr0QrcV55ZP1
QnMi1NZ0LU27E0quIEqlat2gM1+cXB2EyaK4RS61tLinsyg5cNiG99kq4iTnzRFLt+Kz9iGdNLR6
TFDKPGj62cWiF8RWjzyf9Taa8zO1NQWTXVxL2rpYpYXOEZl1Y2mQfWyFgytPqPf7YvR4Mxzn2KxT
Oq7aVlbqX5xzOZBj51c+jjnex/axD63Qd766YCRJW89yFEEngQTa4ACupVIEHBNtPFcf2C+uICgt
JvcEwhA/b7VB7Pc3lMIGJs60Rv8NGCb7tOG4aBIIxPw4uKwgt21JGCUDV+zP/rT8a6YmjLauXDGq
tSy6lb0727ZIhB+73a0csPRJQbxUx3uo9umn4BRAgdlNx1OECELJ34Cz5mU5lcTpD2XmSz0pqWm2
9wfC0qBFg5bQcuFHz0CqDuKj5vUTeIJKjg6BHL1cbsq9PLZa2HYZHohZC9HrfroUzO9ye8xotrHz
y2pqXz6hB/T47lVco20s67xezxB9U/whwgB3/Ub+OnfBnAlBPjbA82dROZX/WY3zPlL6V65pbFG3
/IhUN9T3UcK3e03i4Lb0+ycBKMuImh8OtXyloOg4UeY6pATCVH5Iq54QGn8aK/o5M0Yz4ajAO7aP
9ssWRhRXzwrH8h+HxOKTgcRUDOOjHrA3bIMsjfsn3c5LPaksaUyiDxKZVNnJ7L6kisjkRYP8Un4E
Dgo1lHiAzdnlKEthlXRRBReOHvmrC8Xb2MS7IcsnSsJK+FfOMws7oOMdy42OGXCwN7T+lNfOEY8W
yqZV6UbfpyCqkMz3sJlW5K5i/rpiUXiVvarpxVwAxN8wxGa4KVnxwpMiM+tI/OvU81P/AdgQ9bAf
T+A1zuaCjT2FLAHZF3IpBcnk6aIzGtm+FSP028u/ePmnFrsph6nBkmLyOj5UMSqZGiC1b7veHIyL
+02L3PLUA6vtWHMIpwATfvLP8ui1VZ+cwnC3fPlFRXYcXEtv+AJyLO99+1NpaFNLAK6uAID32hnL
Ek+XbsgriNLLWpgmv5HQNDzoectdhxxjX9QYhkvRbRkyXIQvF3jLYrGC92ElStnCcKDLmUjzupNb
Yop8BbBMHVyEIIQLEx3NgXyoUO97Ui6RAiiDZ8gv7vGOwYdedjNPO/6iZh8516rafeQHsDf+gwjr
4REt3Y6GnSM42YSYeKnb/AZVVFmgFmabN1c+iXA8rupZvleLoAR+uG1kpepfVBNdKpjz90RSgYgT
lwq0tuIbGVGkEe1mt4x3xbaTfjXK830G3VsOBcz2E55na320v/r9S2WUbE59hI+8nCFfjvtVwNEJ
RlXa9GInvFFsNToOMKdG+mLBrtRSXqCKsW5BsFx/RN6mXrEcDVwMPTrW9M8vmwo0+vh2QUZ7u/jN
hVsKCL6SE3izfbQbgpdoiPN1hDnzHEzcs/RHMgGxu0y64nDRmo5lkHhsZzLR9VLdpuuEnjj1d/jw
0rtFlvTbGxoRQN4VeicEcPAc8YRThjXHNNHhmgq8FaxH1iGE2Xtz50J7YBDqIY3BVId5LJv1R6Qd
Ea4k2J0ONkeevbOm8+Ri+tDkLQKjcepYCP9vrbCjm5+9C+KAj/5HRNgvxpfKCkhIQLuVJ6XkkKGm
cmKM1+1orSu4gyoXeQIPfYD/xMOSRBboXPNLwqHMBKVTrlDQNU9Szkn5AlbmlbauXCCSS2Vb5ZBh
OLWhEAX+/wv1zch3xsRCFV4DZLpDsEt9FeGwwZPskzY3PtqttfbtFqkNoWjISMpfQy/e7RxTFkeK
7Q7iA+JMWKLXSDJF9kWvRuIrLpCRdE0MedNY5cUoKZGqvhCf4aHh2ijbx+eXb90eewqra3yreqAq
RcXpZUbBPh8/e0jcCiT1wQHV0SnOuI83Gs/3CE+Yqr2zzsKZs5uX5FyLNmHTAR3h4Ore16FySMLy
R0LeUZI+tIvO+cih6TZGPdV5Hw9cdRTVvTHGFnLxAi6YbzqdI2yYrDTdvR6yIC5Yh+lAjaRwHrtF
Ny8QSdanGrZSQ6lthfJ5cSoYClFJs5bWFceYTGXSyljcIpBPiSZe4SHxpYz6RfeAn8qWwxRJ2Ww2
pb8xJUmkdzoRyA/Azl2MNAs1WCa7rKH9EDTNXSYqz/0WlnpERlT3pfxhnO37dRpLkQLIMLUkq+R+
GN2WXcZ76sSNNkgeH3+DFwCgiECcpL+tGi0a82BxJ/o2fZ59raiDpoQLFrlwtI6+8OTfMsnFpSyh
zxYMyILFZUAPCoLCvomb2cJTP8IB+PAzKdCx0uWzzfVNLmiRBQ9GztKprWHsYnEhrM/sU1iTqRzs
BMKHmlMhLVO1g7t4v4WMVzNSeu9Pxas7SX6iVJ9yOWIbi+yMcG9V8FrKGPV8pxA+b4D40X3ELmDo
yIKiQ3J4dji7zSf/jcfGvgLvv5Cy6ZpBxZa27e1y3jL/JORN3sturNiqVOiuZ9zFCvRfjMADa8e4
Ar/HoIedgqlSzGjFfD3wT8hu5zMSka9CpGwFk63wSvdejMWwDk7WpxZAvvUuzYx3QnNV+Wx9P+XR
fnqOAgwXp7iUjCK464q+VkeTCk7YOuugV3MMS+uXwauStodM7yqM/hPGujVndCqIce8Ro2pEpTMb
LCVpWeMO2YkBR0GzGbxlbfhbZTwbyBkFa/u1XMKWvtcc13CNa2T2Xi8qrkmkAbYhAIpb2m/4Zc0O
B9yEiCGDxsjUoyNN1NP2k8sZuxs50ALBplT7yRVd+cx/wwVNAY0IbWrL3chtW0qPyAHQnuy0cS+z
vF2YRVfX14eunJ57BLw2Wm/tfAja3ncmy3++3qptNoz3IaYohYoi7EE+WpwGjUhhMK/X9CWtvYtn
sk/clD7agL4hd2olcO9lsAsPM6a5ycke7N6BiQadhGgff5E2JuflEBdVeJ5W7euyfSiBOciPdBhG
aCX7bh3Gi0XNiNSZVTvXLxbnU2Nx4BPfAM6M950iIEdzBdyb3uvTJshr/RrqAkswlXN6fKbJnAUu
w/UdT6Fgmc4zJaAjo1YiSWQNLnjTjmdchGvMOAwMVm+gtIUAWCJJLCJdEJhqX7Pl6eM9ucRVHgmp
py8KtnV68yPmDzCLN87bbU4WVCkGzB9rb7UrExDuttkuWBPG8aiQs15AlBzAbPm5FOzpEvC5yj7i
TsHhvNc8ibH0XYsCcLB3JYwdf5cqW0tU4hEzalT6m634eyP5NUBvTqfMu0J49hzsD2lIXB/yG7O/
haYjGYA7vMQ2bMvdSuaKG09P851lWGyXeCNPO6XZixBRmToib57GEutor/lM/dNfQHeD5imCml9e
jMmmuNwzxgNLM9LFkrCxvDKLubU4slIyQnJiud+vzDjOTMdK6kf3pS78/Vat1229Njdscx5gMHNh
oklRnyxoO/BoG7hP6Po6jgZizblb9VuMiikmyM+3YJUliTZuUzn7zE40t5yf3G7M7686mUFp3i/W
rZ/6lzWtd6giNBi2p0bwI3wEb4yiXPgdCyeH6IeMp3Fcw7LCup50p4EGIIoasXhYSzw/QUrURy8u
AJ/YtFPVKs5I4atpzAsVhqeseJOWV5bvQuR7IkuusPAcPaYTMwNsytMPUHxXB9ebDHDwJz4wGsuu
zwFkqBED8snfp1Qz8FximhFR0fDOAk5H7QHm10fSUOcdTNGyRKwV1ay6akE81SYGwuCOcUp7I49n
U4GBcpScOZaylWKZnRkkZfaqU170NRo5E0KLYhlR1+1lwkVCvklyQ+/AdrGQHIBzCeVKKQ4Ba1AX
H8tr2aeceBTPk3h5lJdkN5/ybIkl8oo+GMNrvQ0UDM4lWU+sMubG3orzWHaj+S4nVI9FEfD9zLKs
9hpSUgqK29iUPTaaqyCjaTYmK+0nRXk0hPsYLtImkspOoH9BHuJiG8qR0Kx9eoRP4oyQ+4fhXpwu
jlU8oLVPLpggcr+h4gqpjz6WkqY5usVAClZOHEjVtYAj9fDUqdPCJraPEUq8ubG4cT3Zv4fglHZ2
eG84erY6NhPQOsf0rOKi8TUAZecNVN4bOmz1F/RhJki9gZIjte065ZoSaGScsDsLDroCEoo4bmCK
EdvHIF3uP119gj2I9TNMEZ4N/WGQwYh3JB5Cyhm7998B5tijrDHx5K7u5Ww5CtWwT1Fh/7oQXyPe
zzhlir1rhe6c6rpwWB06z1E7FNjqoaiiXcFlVDhsyyo0OtYP1kEvHW+3dfRKu7aHLqa73HZxpybs
JtVaMgAIRRrgwnWmxpgnubWLmoEYbPHrvjF21d0V6FEfQ/rt6jZhwayQ5zcmJf06uRsbWJ5ylWos
UC8dsc9x4EEkQdNRhIzoO2TQNuNqlhRilwdb4bnYLSzbTpr38azDNnbaWfZDzM+KdEW0fEfDl0p/
nIkEw4h6IRu7kv7BsQ4V9AobEQjwRvyLfThZ6szRqvkE0xn3ChhccsfwDodMFvE7wJv89shDad5B
I5xjiDP+hCknywDdnhUFOnC+pLERoEfnxjd0Qy1x73yo6rQPkL6IcMZ3sXbysNW2uu7GxmA6FRYz
+quvAbdQe9XoProAIQpUAUgpxvY96+6SagtuFnn+Fsz5djPz+b+z1fh14Gv/bN7NjmcmWW0nT4ew
NN7RTEyk8zdLttkzqZkDTZL5sJoHamy3MJDUHrW3c83twdI2TnullR84H1q/dexmCC19ig66LlHF
5Nu3I0OvgH4kK5Uj4IGu8LIjfNLTHJ3G/sVrr/9XCA6nP5ES+EIPEu7Dkka7sThmgw/G3BP/hPCs
MIlr08FoZMdz7G2FqIK3zRmmM5a79Yh7l6rbAyXWyjJNNhMbVKscKpNNk+6oaS4wJoIXTmAIxNbd
3FpGcec8aDHJ16cpF5qlpay+CunYHad/5TIHCsZPfHakEGCwn6qK3CetQsTi0De0Xonky0tJJQKF
Owv9TLzOLExTYxdt17p5K6uRhhNk/59nIaXll/1GYgoM9fMLDMwwPIYYA9F3iyNrUq9wbkAIQ2nd
F1bR7f/MW3YGFEEJe6aWVkynPzCURGW6Evbc54zWQDENWISW/YkOOhJnMF8TmQgwxpTBfwUjz5KM
MU+4DyA4VbjPoGJSpP0VXI5RUNaNQD6GZhHuoeS5hY+mEdtq8K9zE9duGETVAXIqtOnHF27JU0sO
GrWBRXX5OCfm6XqYMcBag8j7/17e1hL64w5b/c7gS4UPznFaUrTsnmRH7+XMep9Zsifl8ZgZ1/ew
ivlu6Yiq7aA49wan2t53WTBGKryziQL3+62huIdK7qFZ7PbigbWuZBOo1Sr2toc6gyNjV+9MgrxT
xt4v/hI6gLY6iF2nj2N5tdKsDaa5J/RBrYrVvo0d/Fj6MOTrhnZ1DSelhsgKP+BK7bmtOSz9LOoi
VozsHdsu2wqxTsHdVkRJuBRtufldO9i8Ce9VGkXu/H9o7m3rEBc5XyWHGWmNeDh0K2LQhmPHCdpc
EsOzaoxjvx5mB/fP4lg75e+B1RI6zRIe8XFAVNC1sC+AnlGVaNvvWdvsYqyAdD6qhOwfX/PmgnDf
56rCmmII/x5ysBnAG0MMVNaoFVmdJ/lSEbHcOqz175eiKXGwqegoQYXS2EFw4KwTy1xhQ0R5NxMM
ZxgiIAzsrB4+AHredVcraET/mYDAkAhfhsMZvhZpjyH3po8904JyiwzRhuThJbsGYNtVoy6IAUw6
VIqgx20wpJRfWzOu8p8gAYvokFMHheMKJgx69HuR1BiyiKLL5cnl3wfpzPlB6anCp/Mfi4S9n2Yq
UE735Oju4eY39KAfMDl31emS/z7Pkapm2HZJd45wOBbtV+n8J7O6k1OYmtSYM1HA37jq/uqA/hb3
DVizhP0TDcOh7G7CGhjPK/6xi+LqSQApDAZEa0neVmXGdhix8Z9KJX3sbXnP4btK3GCxuOOgq909
qD8ulj9MwkGSzCUWDGvlwNAAy0bzFHTjwbtVA0PtmT8pSg2wSS6CsH2Zly/FVICv+Hm+0q43WcvQ
LkwbHBR5UC6Sz2seYpLY/Wxcznzau1iEelpwOC2l1zofs2hODRLcq3o9tWymkdgxe3kHj2VsgYug
CTn5nmPWRCOt2AZcrvTB3E9wIrz9sThw63kKUr5ZZyXo9xypfnUJ4LhbnloMwaudC4xfwXoZTOQ2
8wM8COEw2JCGz25XDmT38CCMZj8H9ge0iCrLCQmGVlbMNjoUt3Vd+jWCQ0irTGA26vezWU/sQ/qr
lInSblLpaQyJqwckvBimlQj+lrWQBOTw0Uva5b0ymmPIFU0hkcr5yXHt5e9GzfnJLh/GZ9AWOgTA
kS3dRttS7Ab2yzyFv8Jjov7mBmqOcIY4p1kqh+NjjzNpFB9DLfi0PpvX1qValPsbBcDIBIq3eIsb
w1FGEyw7nRvwkq92eKG5e+5OHxwN0nCADcjPkS4ru7F55SPDdNe+m+d6Gfmo7lyQ0xrf1JB5OGGj
l0xzbhDOp1Z0rIN7DZWvezVH6px5qfERjed09lGUkJ8LxmDuiE2FrViLu2QpO8G7QnKcB/OvN2y2
M6FHvv31ukrh82jLPMWM0xjvmik2rpAg+o9gZdqxmw5jR0bvOMuaZ9J6I4z/mKUMfCHPEMy1MRqQ
jkL8DsXxgc26ltJfqx4nv8YG9qZnFzNpIlFLFRymBNm5zz427A3f79q4ovgKFbLEvatdnKwY3sb+
Jt8YH0YULYj6wKXme/52+KTZK+E5Zsx9a5gGug9CHfsioigUc3zHWRWjflvmtepamUJ1RDOtxYgI
vJU66O1vkWuBXglPNUXnuQP7lfztTv4yDFDFYXuTL+gELlxTlGFVuSDh29tqfkUhmRzncv37w5Iv
KL6vdMpiGdmMQ6sqXYZdF5NA7jW6KtxsrGiz7SByPXqEjRHiG4erBJOsSUgyoU86EDIlEZCs6b8P
ikgTsaPeRA9u4h8ELBi4RuDGvMA3iGEjhdQR6TwgiIMmQ0j42wiqAfrqnoaognw85dX/p91iZ7JG
IQFDlliqlB/HsfoTuzn74lg5217wBl0ccbWtPiTnJTQrDwJ5c9JD80N6UYAnuIRDvhEXF22g9DHB
0T0MKzT9/Fcq6x4al7kNkxI25na76e/vCBrRHb04ghPSdsmox5Z1udUNTz+Doj3Dls+JCqGvDi5f
uGFvaJyqZwRWSTSdTb9tooeNkeXec3B+8rcMawgcZmARmu+KOGVbrMp8cwjUheqRk9HGB5L9ECDZ
2L/aIxyxYABsdwtOGVXDsw91clQmtM9cIVVbSr4+yIEPKzU+4B97oM2zL7h10QogxacN+FkZNpO8
Ux5VNWQ8IhmUMXgEQjYCu55Ms0yBFhxYyL7Pjuzs69l7q5gBiLKBhR2j3bgD9ZXqwnTHbgptTN+K
c1DLB1xQ1mVfsUdEj1qcReZIC0rAZeMhVkstJbyjCSv7rLov02T3ZoWcQZ4t9bed6tIpXLIYv/7h
pFOdrz+vzoVhf5UugFNhGWOxaOvVX4eiGvycPugEp7deZ3VSAWd4BURbhvZt04YlN8LsCB0vXpaF
XUDWQ31S6IF5oCg8G1n6TU4W/Z79/IO6t/eOWmEiavY09IvyFkf1/55L58/6LLDmoPJQNGF528Ty
xH42BS5IVuwBqrxRg3NfNVR/3e2KUR2+u3888p9J03Qyhd3/QfRVoutnDSzcoEFaZUKenDaxGebz
fkiJhMhmy8JJmvqLD0P0k5VdIEHkA85cYo0UxUJdbZt/ctKpuVJOlGD/quXb1X5dSoZ1MSDqNJw5
vzbR4WtY12o5cCJAbCAjILOQt92l2o2VQLOrwAOhvUs0E2s3Z+uQj6CMe5AYGamnfJjVYJ3a98jj
wt9Uzct6uca9O8u+n2d014j3ni6ZpEzsWfXO/z6SNvDIiZE8IRmNTKjNeyShSP5dMhyqbVMFAcuH
ANhSLJlhWdZDV86CU+4A3LW2QVrmuWrA+quuMMu3NETNZtJZzGNEz7Qv/Iimm00ejPf6Xe5Icr+7
ENAVx/v65trAmd9Gokdgk5RGjXCRASQFnjQgOseGnEdKiJ9wUYrlqlJeWocM2oo+ay6yR2+cPDGy
r5giQlBzEPfwLm5taTPfozN+HZ1o+jlZBQlkHFCuFv0WXDcTlVYGNZf3q3+n/EN2qE9LwWncGVts
9smdmwGg+NZBd2WqVtoP7My1NQmx7oxfC4h2QlZseQRkwOfzWI+ReA0dDpRfsMT97HtLQadS4ioT
i1glQuv65VOOMj19hsRYwFn0cD6TtXYQrgyCj4pyckWuarjUdKMIa5O6KUbLH3jMOD4Z/BaXFrbY
ofmGH1gr7JEN6NNNt5RbsixgsIKXMICE8kaZGWE326d8wnhq8ro9tLfjg/v+SEQdZpN9WcD/XGsL
86HW5ADZ37cQcXcVLdkuopvzz2TNm2BJskxVNqlG9TbZNEOPeA7RlS7qUCYkMtoeBW1073B12A/K
fV5cvrCcLQBX/a/dFagYN1rgEMtkhS/Xrg4p4JR1qYr1IihYVpAnJGqfRcrHPI8N4Auz+FRwJZJ3
Z4/N3HfQ22zCRfRiwYCPQanjNPL7smg+rnAbbIbHHIF82FbxxBoM51NFDcY3E1ILLZCPnccTw2NM
qxnx6t9ddHGdJis6LR+xZk6n6lvQ17UV565NENLJpS8ep8ul4LtFHCVwYxlJC3PYEcBl0rGF5eo0
DRi9GT/05qY8BWNbDOjySkzeXcxsNTElD4BVCWlWonUwkMNjU3rHaYNwdRNpCrG7bh/tPyAUJtnY
yaDnVYT4z+hkmGevCw4Gxx81Hz/CCNfkKxlsC92973dyCGALqyuzOsdA3escy9VsdSjwmaafflrB
Ymvti3kcuRj8awbosBGoEaiRGwGyKE5Ab1dzILAXUvE4+bA4NfApS821lZC/n27sWLFUEQRm6eS3
G/19oVDaW5QfDN1vAfjQoAC4uhU3f9WyyNibC5jkvUmNYZDFRKnzX9GdojeYiZMw7eIg6i0dl0Ya
LdTesAiHzNaA/UQCdz2zyXnDActDmr0cyNbCth9qFxecejnlfhelUBsHShoU6iVvcNq8BL1VZ9BR
qD2lexaOtjM4ZMSaH65LCsVAMrXbJ6c+fsHzbGLwSPxqnmnJGY7T1Vc9dCOCb+QUTO79n8RErlVC
CjN46+O6DprJnAMqgmSFf/zphkcisBgOBBWdNWX9fMnA0S5pI4Q513DcPk2KbcftdQPKl2WtnTyF
zsgR2ocweMKWpOFowkRKjDOlFhnFQ8H3867VA9sSC7Zv9n/VrJzPM6o65+eFrn12n46BNJ21PCfd
Rwe2XHhKMdeYLRezAKPI8N5JVy7vlIN1m7iLMKEl1Ei+/xoYOqB2d9XdwENpOt7G6EEogdRFd7/l
x4Grly9aHoze1i/bpyjHmnPmlp58sqRNiFc8lefGeympWifDtASYg5f77P1BzUw6Q+tnZAGY3Ny0
GDIBTqWMJZfDJrg0GUwJ7MKGMpBsdGLgPe8Q5rTizibddhBM1tLLrUMygGpzhEmwyXOeNWhQTViA
0EQzYkOuJwckLRTnsWOvZtJZLm1VJByLk0nNtwhEcR/bZcmoxzc4kECR7gdQYG6iY+DdyqaUYXZF
m3drEQU+c7kNeWSWh5sTtuB0NKlyTFsCAxQvn0aB+t2tS7GwcqcSmg39T93Rokmgd39AYLcNy62I
+BEBlyWOOaIp9QqwW0sCNeOn0ph8TKOQivofghTkn3eQ8WY+ULaW2ttKikMni9p2lgq75fcbfFli
L2ajkphb2+Ex5bngDNiVM4JU3ROUvlKBCbiADmfppHWdsGm/FYbHpWDzqs1MiGSX7F/49LLKLeb5
i8BtkgSfru9Fai7suOocQ2R+WosMsbxSUidSOIXqDMQQpb6QOYxdte7/RfrSwwCXvf3kRotazjhL
7E4OcpgdfNqmzfw2gx59o3iWub5+95AXS4bvGNOldwevVPN164MRnnfzeuxIPks/GRiRGdYD3cHG
CdRqOrt/5XP081GbSDZ6ssqudf2wEdvP8zlxvakzekKiGEd9Vdd+7xfgXqThj3kGijDiC5U8P82A
EcWw81dndOv3TNauXje2ApXniyYiiQz4iNpyEL0ahPGx94cPJ1C9OhWUFMEC2i7DQhUs1ls+k/0g
MXlhV/FIv5F5l+bn9GnPjd9Kx4GKOEl1Qib1MehRFfvnAUDDGYJZSgpYPxVKPM3rjHwnZgulAyUL
68RSVnmWBD4LQgLqUMFvhFdoT74B/iY52wBr8GXQidCif9kRVvY7iPdz6VRgeTkUqkm7bj4bO1SR
+OVWx5UXwDKc6j5tt7i+Kn1YUAbd05Noyq8uaBL2NdqVB76eXJZAcTZFypv0k/6nvm+QF6bin2+3
o1OHxlTwQO78BnTWRyuDmZLLHGY+bkIDZiHKKyWK6ICzXfATPVv6Ff/zy6JEjnbS70/FVsP4Z8UH
7RrRmR4ncqJA2FWQ+g+8i2BAdlDXELUAPM38gt5rlLyu0pr6mG3pDeqPZ33mZjyZyey3Trg7J0t6
saLjB07V4CLupr3RVTVBVmYdm13hObGXC7deldOJpcfvbOjD2dJja4vLZBgXB2z9/uW1jCBn99Oc
SsGF0l6IOM/TlQ4pjLBpxY2MBvdpiWpuyanY1dGiI/84tHqi0coiLt9cZHAgcbOamCJ3fvRFJ4oH
5UcfJ/nNPxlZUR8AwcqSAQD6D4z0wad0hSitbYyF+xhV7xgbgNKoXKD+9HMvU2y1ipYa/Ih124cL
dtXG7kTj0d97xqzL5if2NExMo7Z5k8juNwP+dvsTV4vrXSqDMdZKfWaKy2XcrrJA8EF/nv8vTON4
D2cNAFv3geKD0EpiOxPEZmGL7XQyBjFtcHZdqU0aPvMwF3Zq9WQ3nQjARKxNh49Nt0lUsEFHFRox
eR5SM2ekitRDs09eFHShOkYNlVkR/A1K0IN1dXB2o2PJDXoJIpIQfWMP4KrPY2/h2KTPK7fbeEu6
rWykW3+L0x3a6Flb8rskk205i6FR3IXzSX+HIfGpjUfkaxvjJkwYIGlowwwrs9QY63rh8P1p8U8X
rgqDN40hRkADoV2zbJjnswQ2qAIAV90lw/6pM30v23r/ZmFG9JLAviuryQWrezN8rmMzTGf6ceJc
d+j9pXVwtNXT78A+s1XiK+ucbVOm69d+RDLsW4SXhxBHjPL6QVmHVQK8FKAeLfahg7VcfcL/z762
040DHNPajNKBEfHzME0f/sDpICEdSzDBvh9ktiF8WSbL3LzXFj+n8j2r9kPUvKiY8b1vDxJObPXX
ErxH7tFgM7LgSIRb6bpuZ0CIIy98K6v/L4vsvXwCXMU/vzPiwo4SzftA+Rd7a4TliuQIY6ilkJfj
e66TTvskqLVtbLHSD63WUqm+NBWrZxDZv+NjJ2cpLf9VwlnUuWyb1KF9X61OeKwICV5MWkScikTM
Xt3vRwuoGmSmruB9wGhdzNWLVlmQQ7crow7opCKrwaqHiYGirUxb2DQpMghZk/XiodWk90dZEhvr
JUyalRtNzJ4kojeFCiU8FoYudZOQX7gII6o4Kb01Whs3lDJvfhWXbTD9eKz4LqfBGgbMvOJSLNoy
RDScv9QZQ75Jznx9yjr2UpuytjXvCJOzKFP/I/LC74ZidzvuwpJbM2GQ2P1AT+yIkAwXrMHqZRVL
eBwwqAC9PWYacaL4zgXZJXEpRKqItjG+cyV/calvnv9Egh8AoH8qHQ1b8JvtMG3TbN/A4tHJkE73
aotjUj5I5DN5RMsDwKWNQqX7gqO981keJOygUthFUaK6OeCvk0KPaIH9Wx6bY51AHD64Z+po3XrZ
/ZHTeLhImfxlU4OzjplWmvsKbzdZlgLwI7LAAFdxpBCcuvrlDN9q8jDR+M0LTJwpGl1j9p5XJtn5
RTvG6/TW4aAnc8Pbo6k1R9YcAZ7tUmLbFA9tjftvrHEiqRtH+b3RLZVrTK08eY1UyHsXSFwuIAwi
10KqUbiXe1+1xtNZFg3lpcEU8sEaXliTp/5tG8Ebnqv5/lEihIQUpYRVH5VgpgTxXV5/siwWJ7Ey
Tjimy/OcZUqdFF7vRfqQ3jSgVK21yrGkNE+Vh3I30wvOIYU1x7xx7Z3kgp1hqOA7zxIqerf2m+7A
8CpajWtWxd0aUKUAPH1f5Dt3sOPsG1xVjZdFVTe2ZzO3DPP4ppSpYtN6xAm6gSY/mJbv1MXVsrgg
TCtVjb7C4UFzu7VohLmBudr1CrtGqWJs40JoajPLHXsKs8EV0h2PvRPOX86graPN+dAQX1M1iK6r
OZG+eNqlHvROrXh8CiHkNvRgb0gkfIdKaFarlu/UXEpMPhj40FUk7R9ARNp/OZIrwtL9hkrOkZyT
fHE3XiLrAyr7rVJ36V/9Q2uWuqAwpssK/2Y3qfKs1mJXTVOSj6Ea1/HJylzsF9DSUbQf1syAxfij
x8jd8fYMgMgUb7gCZCKe4U7de+JSNaYIH8Hb/zSm60oOjN6JEX7oi7N1ziyWGDhv2caQqMpnRZK9
q4LKQSrvYyagIfNkt4EFifs5iu4NVUgC8N+0DPhwIiQ7AeZXTQ54B36V0CYll8X40zcj9K16bFYA
eyQSI7GyVSGoTeNV9VP+TNiqCCndsXfeQ9l6mOvaASTS1B26hRefQW9ZVmTM7FHiys6n6Zy2H/PF
OeYoFkpau8qjc15Kx38XT9Sgshn7qBhRZh8SdKVDT51Eem7i0LOxSAKbLhC+9eEk1SlRr1zQQAij
0zSsMFAh7Y8FxU85fRSdt2U3QBVDyWQ864CfOR+dC814t4nun4Cax+EYxplCFRPIEXLE4ojJdjvC
SV7TiSiu3JaQ5fl8Db9FPt7xHMoMY3MO32BlFP/HkuQw1YZoeEVLDai7VxZ3CkmUqPcbQ8W97TdH
WymCId7CI1HiUn4rpz7h9y3xZut/Yc2s/rDkNXd2vbvL1hCu1SdZ04rn24FvdmdEnamzvM3reIeQ
1npukUVZj4x0tqUr2KoNRpbjuJINIZZrObheI/qJ9Ns3SymW5qIAZWMN6bOBzrstK/b1pSN+Bc44
A63xNcpCYf/JN5VmZ5dZIWLGeEoNG+ddebKi4BrWT/A7FQTh5VI60IDC5449Ydap33Q8CA4Lowkk
EdgF0jL209fV1iMsA4JX3suwmBBz38scUO/5xYvL7CcI68VJHQYo+klCiA9IoCQuCgkk/hh72fHs
IUxY04j6rl2vMSKLbRDT/8CTL0h2QszKJkzWLlsIrTHUYpa9zAx/tOEhzmwuB2VSvvvql7MKhIa2
7LbyJKRyl+JqeCA16q9DvGXYnAOIDnj5O3afadBmO7IzvmsD51HWt7BRHbn65Dboen9jA32XYog1
rzNWOo8yUdCasCMNnoRjbiz3Bmh3r97sfrAyhq262ZTSRObNAZAOc0HR3K6ltQu6fKAlXnZBerRb
jjQGyAmBTibdrai1n83pRG37CRH4oR17J0da0TAiLe76dkCpGScrj4O0LChyeu9J/+MCVMZQQbR7
cl7rsmTcsDYqfL4K5/K73pzfktaAlvdCKcRTkkvjNZo4mb3ja6y439Xb6IQ246aXDCaK9Hf+kB3k
OcZkNu3eKF24liPhrhB7SFQ06ilcE0uGj5x6LbxdylE7kgIrKnTMrP1d4PcxP8mGRG4T990nq4hq
r8LjYdtzFdv7MqLMmZ667wd+p3OvijGjRW5b9ynoV4bmsH5ZLX72OCPpHUTfKwkdJakBO+mcz4ki
AfTM+vAC14KFR4QXIZ9Y91VoB4qH8Dxxicls190AvwrPhqbi2Kgr4mtwu3tR1LxyTnPgZ8xkJm3g
1KL5ZNefb+T6Xsu/MrWOm4LJ5na9QFonHv365/UgJQtIdmyDN9csoIIB/QRJQotfFc99+Oz/0n9p
fYI4xB2+y7PD6LaXYlnmovNAeFmqpzO3VWO2tUm0Z0fWRmNZSuYTquc9XZrkHiJ8+Uz5hnEN0Xup
Pddb0qyVU3PVl01c7YQ6zZcFdirDf+B0VaJytHrub9BLW6wU4fbghD/4bUpd75RoBVmlTP7/1oVy
gJLYoL2m7wW/qXuiA5rP6vynJMS7OFJIBuo13FYyFmvnu8gKh70bhiemc0mmDbKQ0xnmZ2t1xYY9
nUHqg0kD2WDyhDuhmHb/bYHd3YlZet//+7LdvJdWPMv2BVV5NwKibkZbmlAxgAmGlwH8tKi9H2dX
ucCFoyr6xtjIAkuCkEwxE8S9q9GbWveRQLaXUNhB4DEd5m8qhjW8uXpDCg+apndrV9idXZbfEMuo
i0NFSd97PO/MEbSDnlpS0rdSBbaCkIFQh5f5NFM5urBE9ryvvuyWBSevauA+d6+morWpZI7w+yQM
GJ+00CTBirnKnPpqzH9Ed2suPGFRND4HlvqR557twWb+WlPLlcse1NVSgo3fScBdexl/Lw+jbaQF
rEBb8p79ZfBVSCneMh5vC2O04lXtMy4ruCSygqGKWLw+rdBxtkSe7/7IJ0ZX1iX+k85ZMqZ3R2oK
UF3D5MeIp4qu/i5GHjusjh+7BTfcXRzIZrGvZ9NJG4kRLbO6zAFL3C/pJwF8fgW2oCqPt2sm2wy3
TPPriX2W3E8nW0K3iG4kRpkkM/RCthZSWIfUnS7jfrtjZpvhyOaFQo9RPlGNf+x7WhaX/3DgX5Wv
gQkF1ngxDp5y0F1vBfXZRbiRIBMZB9GQGLYs/WMJlihY/iHtbTlEgA9+U714B1NnGf6jF28Nwrz0
29lBWNZDFJp7C8e2c87+PS92dQNF1+fOqgWsHnfvtqGx6WJIVxzCsuFkpM+f33v6nrtv7vMyY3tC
URHEr/RYVpr3feM3EeXnAUXOg2fdH71pPV2cyxwHHUab8LTEHhL3a1XB1AVx+4+U38Iah4/isFdV
hzOpEzVOLEElghxURHZddau79l1CwFi27p4JyW1eK8hMaaFhJtOYrNW0b8WYs85FXw+widoNOTvD
RAV0N65dhaEpEW2SxDrwlwyxUUMP+5YqzE/BHdnosa80C0gEwqp3FMNsahl+SzsuCvH44VAbNm4U
+qXGCWoZ2uysM3OD5TzuRZMisSPL/uGb/IUmRq6AIPR6f76+YBxKoUJLoAcUmGOgfjcmtBtFmaxE
+gE0rsL51GskaK9dH4aMgGW6qI6jhMG+mZaAgdsFIaku4+FNP9c21F/DVjLU+aPwZooI5PNgfNuX
Irtr2S42s4W6j03neWGnkP+97a8BapBJ8ZwZQ/nc9E5ZoZ+0rTFA1skyF/JCvEbHqow9Kut4SDBo
7sN4KmZpuhSCAciz6D0iJucLKBRmOO2siWVPldzY3G7w4MASg1Y6UQ8jXUgqFrYE1uW0wjyEpwEF
d1AE2zZ68HAG9jsNlMCHlEIa1oi4vluao5UPbSZjk5s5YqrxP//Ei3p1hhcRQ1KPXjpQCONvaUFU
x+Ku/R6kHwIXfCFJd13H4gT8Z5b5jptrvGSKRpeWukFCYfWtsQBG3OP4QBRQloRpy7NGgHBgHURk
o5Mu1jbS08wmIyu72mW3rn/CjQaniK67vV7ZYpCfjtX0ffaujomiz9tx5YEvvZ3uzeCEQ94tJky+
4F3el7us1saxojQ9U4Jo6G7910jfXnm4JjXoMWysN8zPzSLi0L+NrCfLi7EvUEBD5ysw7CaUB8xp
EZfLawvoZEGpJEziOD5qpruW6VPlIvyfu6mSOC8FIqFbOc06UZHLK8zdBcNw1aZmzJ7xn9Sz9VMD
+mjhxo3azuRYZKA6RVM09f5TFBkO0P7R4CKKAamEG9pGUvXgwXAmG6ijFwaxVPKvSBW1+jZYV7BP
ylRyWnAKp6mMGF4jGrgRZXt24DWC4i/PeQ+70TOCY3ki9nn+jV8aqpsEmusm3TWNoQW1yxqxwR11
ohGWyuNs9Zy6/cjVKXdbZIKKnUq/Hd9LnEbwpbVM5SCU5f7TpDDqOKlF/K5/JNf7SsH4AEERh/hH
0M43yyJoKU3nraCwQeVch5ZgrJGrWUr9+fJIlN7iwj/qGC/J6aDN/fgIBqHdHlW4jiKhL7P8LPhV
4qVdd5i8fqO5z5qpVfFBcYftdkd5Ol59/9kdz5Gb970yG86R5zP5EjRV0QrJNV6pbMoUcjS7VySA
8N3eU0lE+CwoujIaZOwlXP5h+9FktVuDwsaXov93yfkJ6cx6BQMPNJ92nQ/gjNBhKyMhtKryp7Ae
HoeoAr6/64bT4BBU+9Ae8si1yeTs+9e6ByE4vm9bPfwc99nHnXTnl7bBfTvwnQlUgqEKmELTqB7I
tck3XXvXHR3hkxDHUYU1QPWjBKtHNL/WiUGaZxNHVF1swNEmpBDFZM3s69r0c9Pjl0AaOF6TfM57
+mpe4SBKUIVcDNgeKmtGKYrR9DSb43ERLv5WFXnwVdmsbETd+L8OmKr7oY/fNcBukSD/PW7WYLc8
nObk0JRqa9ZdCUg5cwiBseQAIxboClGkb5oE3bQ7ivedS4ZXCWbhQBltmL6uDgf2QiXPK2MJOvGL
TRWnCd3GIIW5QMxtALUCM5Sl0rg76K3C1Fun+3JU0Y8AYh8JqYTy9Uwk56NfGwCU1abFzikMgTqs
o+bWYtgRLawVT5f69rkzoAOUlvVRsHPY5xSOYvi+PkX9TVw08WSxN7xhIpOMFQHB+0l0YpoZjXuv
rWb7JyZ71MGgPNvjHHXFbg1jIyKGG+bC6e0wjgxd1FOU4xG5KYdA9zxbgIheeBJZPyV4TTZ9FsHJ
j3oRGGa7e+nE45MXb8Sx1JZCbBYfMQI3gh69pIEwqpUkUPzPLAPXsdvuye+7TVYWELUdWL9NVRLa
jP49p07VcxNnGqNsuCJ9hn3w3f2KTH9V2Na+49ZiskOOjkbR+1R1rc2/n9hR5/OWwWhqmi4RLFYh
g9pnvptWup5XwqI48iupB951Y+mtmhsYBZasq3EOCp51mg1x5u/lhwvZJpfrOqE5biEYOn7qaHZ+
XrR1k9bAN5aoHGWZnMt0c8mPstdY9Ps5Me47Q+MeP+0KF6uAGOW+7mw0glyFwgJADciqXwWSXZNq
px0iaafNI58oiyGqXVwacLBaYUg3FCCIgd2RjgSQHWkSiG8lXaln1/z3tjh2/Qyyv0JSLzFiVEJp
UOucofTt0oW26tENrVkg2r3UnYlzmBr067QjJ0BDTlXpT+vG8FphCh0W++WfiusjV4M2WrYFDXqR
74hU5QOpeJsdjgz3Mf2RNPGy8S/M3VKy6FqiYj4Emo/dA4lYT0ixkzW9yLCpqJ2jdNB8QWndlweN
vYDhHaQBp/eXWXxNoxVKv+c8mjCpWiBVcHlBlOSlJZn9bokI6S1nRlHB6d1yjaA+n+530Yt0MKug
EyEukeSjR6tFpnMBDfcCAL6cHgu6Nm3e1wGvK3nBZXtOXmXHM7ukucEV2TJSl39G5kXVRPDRage5
ijac2s12QDG9oKmE/94GZpuSFVvct2zCCaMA0f2wPo61OI4qEqCCBEutPtQqv36BQJaPfinuvsYn
VF9v9pXqrEvx7NCjKpm6zUXmws7AzOAmBifV+5GxrUsU1FBGl65UGAOi0+xzo2ngZpjoJPab0npn
e4XRqJfRBQuzTmxHMx57vmA1pCKCDCvw+Ijq+v0sdBo/dQJ3FCJrsSUN0xZWVKFJZ6nwkOaiywOX
z3iTFC7lUZ1wRElraoB279KEQ/kOFb0zy/gFJ3q0F/LDcnve1bzAAUJTyvP+NsYYWPrbLUd9RTPa
qLjaJ6H95RZuGc24kWtbwyzItEUDFsBhNcIeFCsfEP1iehpJrtR6vSgb9AJANyP4X8zFjeITnUX4
wJup6IWYjICtAyYDwRJaF+sCOmpUdg+ZOIycV2f5LR7oCsPEhj1uScWX1x8isMbOGNSlGL0iH3Xo
elHfR/sHnK/uvbVz2jm4kGR9tkZh3lNM089RC9TUAEY95Zb83H7eBk+0oamsS+0SD4hdF5JNr1Ri
eQq+mp2HE2RHLka1RnOYA7PNUnNKaduCVfhxfbk1sd02wq3eWplMXUF/tTslq9IlwRibRKp+cO6k
gP5c5IjmgpoUP4ouEZdkeehu8bKVRO8QfFIxSTw3pU9ue994A49KsWy+oiq+R7YjXlb4a8EuneP2
HWP77JdvcIM45jQE/8MZ795mZTEBJQDQNjEpKh1QHZqcZTHf75I1zauJXAePDxrU2LaawEcOCyr9
yfsntS89j46QfTakkscgvCjPfpyimUxWrKZVxXCpQED/osvyHN4/I75XXf/lVEd5k7rNVIMFn72y
dJg9fvG5XNNBxDoa0WjDs4+YYpN7exg2AHlJ1FQ8FTobutEutxwHP2p1HCWsvlwfxe2Bu1m3gwJ9
t+XdBNp3zq5HWK2TMsp6KeFR+eJJEAQm/59MnevS3oUlh9sNXJSBv5v82GAx9bz34q59yErz8St/
GbBP1T5mpKPTyqLkrBvAVIwHNfKwAArmsDNqt40YRCkqCj9fn/YDD9dRIj2AoY9sTq8gL6Y9dwOt
wMHmaljW3P+6dSg7HAr80N8+4879AzKw8caGcAL2rmSUhG3FZjsLZV2If1scdq0S63WLNkM41rIq
Lb2UZ76/iC+7FZYWaUrLc5Lsuhkya4j3vN+sQXnmwPmycLmQvU6soUP2fNoyIr4QOT3IiSS4nPLM
LpNJQwj/CQ+stocLbMKAKeYIYQehDA1r9ncnKE6ULZSAgrnefkIJFCfkd7bbd0k98ofbvusVonHD
f5qy5VOeCeY1HSzfX21wSRziSpg25MQOcWJf3Kd4MYw8DpD1UFo4Tq9bjCNp7uLfvv1aA+dgvTgn
Sjoi/jGSTmKowOj8TiJtM8HHkv9kg4Utq/JItdtTU2Vc2yrBdVIyM5edxYctIXApMArGz8u/juzG
w8kND+EpBM6vHs0UxYyEV//ngj8HfG4zx9KXggxJh6N2bgwXYd0yVHSnN2queMcjgMAm8ojmyjOf
KoCraI+R5PZktcVxKpJsuxXV6RJ+osSiG9zvYl4hJcUmsQT1cAci3MCi044LhZjOAuKAeO8l72HP
OXzcorBS+0u60ZhPKvILVknuEUxo2EruqzUWLxVKMMzsVielGgFhyiDvmghDMc4LvXscV2CWx1xW
2sCwXGBKac4/8/Jb9tf0cLDhDk/PF1amEEB7G8ythkCZ7D5+Ko9r/W4z/nmiehIpwhjz0eTjY6QP
aiYhfmzUomFTw2aWXh8XCD8Ao+UpOOchS4nLQU2bGL07L7MTkU/5radZIGacluCqI9Bued9ODYCQ
3zhWjdL8VQc4VN8wKqxo+vNNe6KIDR6MPdNq9dnQmFI7iBwaHdAHcbEy8HOtwwr8herjraPSpPy8
dD/qLOmRJCeViz5Xzmk9IILcFWL9CVN+5LxBLkHds4/gjiXC/NOuxXJuCJAp+FnjLiJoTTypP48Z
XikY6ElBffe6MyHvZGSYvXRGmfZ28pi21ErNdI6EqBFOR0s88nRR/EfjSafqCE8pqKPvipXTGuL/
pqV74r58eTd33G60Lp5hfna5/7yGCCCWZmMpAX1fVx+D2YAFH0clxXCQ77UMr8M4jXIDoy5oosDv
FVJP15V2kGYSerh+PD6gKwkci1pfC/T9/UgPpsL5+xGwlh7a+2nMjJM/BUaHq6qSVJdJFOnaasLO
qcb1JTmCdvM0JgSNE/iNl4pXAziaXQX/YSv/J7QaJlaucYM8wY/5Ip2NhvP/fo6O/EjsbQWrK2oM
0si98iXyoHU7b8T74ExmLQ7J6kChmsvuvbSfJNhh94SCg/8DcyRsHkZwv4S3eWhX1jddYdezEKzc
2wjIraUq97ZeZcu+xqW9KQ2g01x5yOLZO+iKesrcN1s2rK3sy6bHew0Uei+jb+LnMWSsrqhWQ8qQ
oxTxGhsanQ4AiUWmU2B/rNEjnXeyv18k10+nhOJQUF+Zjth2DJSTvVLmAYgesGvKeiF/vqasu0E1
NOPrJBzf1xNPvr/7GDnYNTujdarKCCgfUCHxV9vkrLK+czP/3j9CdkgxvMiwTArLDI1HSBq9CjqZ
3K/vsT3HZJj8Yoq1Y1jO+sDydkzB/VluAGTUChqGBnLt+K69uTfYDCkETnDm2QUwgUFxAERi6Ihw
oveb9d2N86H6acwI1pHWOgMAz+K2Qx6xpeXCXurbRJh9y5IBWUGCzcHLIRMYypkACXykTPu9LAcg
TdcCrqawnry/3dez/m+3UPO0mydx9Q5RWQOJ7nvsl2ZvP5UjGZ8e8gjXG9Er3MYtaKuABqeuzcah
biIRMHmsRqKhYK149LwOaIV997sbovvaQ4bbbQomjETUrUctlp2CQiPLH8nlqjKh05s+AYKDLCYA
KiLFl7vg+6W7meaFoKoQkZF8cs3IrWkMqI2gUshSxazlgrB9XWA0Y7bZwU6pHKHglibmZK5oDKl0
U5OtRu29IRB/9qrwzMQsE5bnb0qsylITVgW3iMemmjzIctvT3Gh6Z3ur/+hPVnV0EFrrBAMMRvQ8
NoxqvXQ5QID638kDfFAD6hAh5YUBUkzUq2HHqFYqhFVoYwwfhs5wCElxc3pV/7Zv6uY/V0pPSZyj
jarxH6/055t6DSCqzg+p5yVz3otgrpL9kFxmXXS5LKBJ0oPbJOTbb+xCA5KlLofprqh9oX0OQTcb
NDfNbqbgRICN8pakCNnszTrjoIz/8Lcd/p3AshYN4DXrUEQeKYrB0LEHjUZF55/foPKUfhVKwmur
zX+FuJlrkS/7SKMemgbKINxKb3u3x7z34XsJrdt5b5r8GBMtQv3yTiiC2rLG560jpP0OSke1H/XF
yj/PkkQVAAkiy8GrrxU4vxQaSMiUFL0/leLiFgXvlzI77UpXVgxuuSHOZdD/tZxq47CTwsHPEFyq
DCJ5PAO17SA1OOOATFCluLQMx4pKEM1NTrVpADEHnlOsf+XatcXdbQa4XjnDPn/Yn/FvkzKXcdNH
Zke7Ugwpp06baAxXxJvEqeNYDY8COTMPfNCqxqvU95qhOlf/ML4dKUarI4Txs+VVIfmHtONRWdpE
Ug5a9J5xx25L/EDlaL0KGiPsb1CcUTbJrFuCIwUFVxfVdQnSrj4Xh+9o0uipB5aSlL0Gnfb8UDAK
6gMxWMY9b9SdrQ5TetzkQr3GhHAAZKIZ9hcEYy5DpBoAlquIP8b8r2mnS5xkfUDguYLF1VkbDEEF
zsc6b9uXky7qphs0C8O+iR97Ofxns4sPhc+RtJ4j6uUNArvf99hZo/CnOPIwMTaCgZNZPj9U8j+8
b15QxCC3/Z+KkFNJWRmzFWFfQSAI6tZrtzXHqDxEw7924TvGx9rrnay21aGHtDlYumMcIRmPs43g
t19ofzL6j2vgT1QxKceWRNaUK6R1ukOFBmy+Z6lHxbsfBOGg+SLKFW+l+C+1rkoguD+AS0ITnORd
i08fr0AGBdgipfmHdT/lOpk9v7n/U9LM/GpJ2+OWPcDESdw4BNEBl8F/OyAc56xEY0CWBITyNSJC
URFO5bqQj/APaX7focxYBJ/epVDk2AruLw2WU+s4ehEznlKW0rcJhSKY4oZy39ALwkE35Tq1z6k8
twtIv/pjecTsp38mquAmv8vpzLmtR07tiyzrYvrHP61xoeaHkI77TXG8JOSVDhwFm+67zaDvCTfG
1Y7YFx7XqJABtpkp5ZMi1FJMuQ9A1c7oXPMl0NiWdyey+LoEdIkwBgwM844gQTzTDf38OcZrOaSF
aFlShi8yQfnpxZ0BzePO+Kh76rJoKrzv4EFAhRI60kFecHSobIvGmhyVDV9FZmk3X6Gy90BjWQaR
Js1qsWpytJTGh0DdiTlNy8bqTn0zef1XM4fvVCL22GmlrchsqCvnm5K40V+luTsuGvYvGD9th7ud
X7kUuBMywx+GPKl1rU/w23GeWslKVL1Rcn7Xq+TpsqEw5v2L/o403b7piAhPqVvEqS5sCEmqf/8d
O9o3jDFihLi01257W894MnTFWcZSPi/aBDOqCq3bkrAHUD0EnCYqQQryb7f1ltoWUZWGkDI8MYhd
hLOMFmUt+C61Lq6Vjhs/FGmt6MZfUeIcYo69CtXUXLteGWctYTmnRhsNcugOcDUxpen3r2xZG5LW
MrQ1yPTbfU6s7/VJl3pWA+DuaTCdZR6CfwkRensbMRkdNkSVrd4kAEhIl7x195CaFxM8O0kCNmVu
NlCS42ybr2t1uvENZOT+bUEfOTI21XEpOGxpNbth61WQMcE8IHjiKQ7nJEptJmgiI/mMLCvlxgVr
+FdUYumDf2hYL/cdxoGp1x1cwui0YPt2YCXlP7KZudRE0rzeTCfhbesIBDiFcx+xhok/oLfBsDeA
c/PRiqYM5PxXdK1ixEwyl3RQvnQsn/eaBPDp1zCzVuc2M/oeJpDMDSglj3nClxQ5+3G5tHuxQ9B+
8h/jkB9vdngYQRToRH3LUUqC6DtgF3n4eF26plc6pYrYosHvFNR24IUzrCDResLbb92x4w6a76ii
hHD2qVRm2TCOlpQJ+mB+5alUC55GAW+W6CHhllDIBdqdml1AiFaY5hIFXHa3Z9YKrs9CHjvbq+aL
kGefHeDqaYA3flnZXCoNl458iNYEjZ0eb/5QcavwLC6C/cr0y0fHhSqYCfVwOQ6Ci67jqHPfARIw
aetpXxGiXydyFBFeS3WkUcZds4FD8rb2QoO2ccgDSkDKjqT6vhN3UVdtB+IGkPobFOEjtKjh8GII
gSPquEAYOLpZSGKQo3c+ohDLKewA6Yb1nvth4mS6A9cp9/ch847YHNYGYNsOE8ojqD/Q0Kz6k6en
PrVT+reILjIPV1sGt3iIy2SYM+roRW/aqljyGf5k3xlCPwvn4q4Ti+fOKyAcNz+NphP2wVQmgSUJ
E30dgtV/TTulT2XRUZcW9cjXHA7SBYtXdQ49xt5RHgiwXQ8mrf9noA+0P0qnnY7JoJznSUd2sQcg
SOZdG2ts49ewmYTBJxSZlfPjZ9Ac1L6UHTplk3e1f8Z3q6l5hah6VuTzo4QRbrRPHXQ8DyXGq6DP
18LFb9rXk/mbBVJWErmuRd222+8g8M8KDpm9H+FnA+5WQF919iF6lVbXv6Qcd4bIJNfgog4gDjux
dMl+gTeyxu4RwGs5dQ2jx8T2+ibsbEtvbw24901yPQk77hsBB1PQt4UT/mtxSNPoyELL5GLJdlFu
EvMO1dJyOFZNwY8VjZRcvS2Zd3/AkLDvO8Cky+qVsj7NclN/cKPg9d0+FfbR3FqX3rPoRE4EQgBm
y4GJhGEU0R9BWZgPCtkILEZkeYskbUya0roi9ESBLW0sZYtvJFMZE/xSB0qz91En4c7m5+sf9+1L
TXO9+b9Fx6ghmdC1hhgH7aoKwC6+qDl/4Bv5/Qw2qvYvFzd/43OO36mQs/cLu21C5Uhkg+MeRX4g
hBZ5+5+FfUtyjrAeY2Kz9HHfzogrbD6pfR5RANVmnc3ROcCs/+HziRrI+h4ULD9jGPS4EZcV01Ud
1wMEY2FNU/PRyrJpM6mcJnSby+EtHufP9NgUuOBgHz2n2sYYU3K7ZUxd/0OAeIwLR++ci8SlPUfe
rx0sHcHjqmF3k+xl7jHng7N3hA1TopHviowPhjhNMeq7yEJL76BKn2X1wBX6GyftsFpSPi59D16Q
ecwCL1drLd3oNhJRtvCJthmhF81qxWG2I85JI4QyCVRsJZlZWfpvuONhoDGugtBIFM3dmGEIE4et
lVb+bZWTwccJ1uq1jxSX44n1xY322w5cA9DwFe3bJIodkIrI7zqqm3Z9Hk541TZ9T26c8uQ+GChu
vqt49z1qUxV9vey+z7yapHigpXZ3qNnPCPHs1FXA2gOL0iFOpecgS3HnmvcVCdSrGFOHI4JiZhYw
Py6kaRXBZcvMNUGzAbRoXHi1iLKUB3GX+e8OlclnJFhKLFPicz2FXEIWutobs7Q4qEAan6vv+g4m
+njJEQUEkInZNiT3JMb/4jNtZtmKeMAdTqtTJjabn4+ANJgf9U0uwSWFUlLhIkAJL6w20IwzYzRO
naxXZMbGSCRUECHAQW7ee4JBOQbgYJoTGjAmGfM/1dVcuO/GNVjp+dA/09iUnjTuUx+uyO5MiOss
zAc7Q00wfkkF6IkHjzQmfXpNd8OBJjHdOp6D/4Tgism85RcBg9AmxDcyvNofH96/p6hHO2qwGvC9
2rmohV0hhvTtBsIBOTekky0lWeFjCpzklzKqINKWSSjkO/6lpUsyDkujSdkx7DoWjHMXVZjs4PO9
Rp6UVpIsU72rD5v9bbe7NiQ450zLW44tNZCO8fN4xdiBYygbKIEFopjCAG3ELSs8mGgW8Kbco9qc
L2Ab81CsI2A58XlAUm6SNwj/MBBLbkmfeaMTHG3lvZ1aS7EWVz+FBXfodTRoaM6J/1yYLVm2m70w
pgHgMSmNAILG/e0ec+bPjQq/SbUSakYRmLAwp9vvCQSrXxGBGhh+En0wnKKXoo/oDViE6qbTvjh3
u/eTqyuMguM2AnuV6N742TtJhOs3fsg4lkAOPY9C9SGFqP8VVN1JnnS47NxehrRzr0o2HLdjYfAz
bLn8ukp2JCvQ/ejyKGCur4smyxS8GmJccPVjN8ZMVsr+hu7pGielKhkAhFJXM9aROhBCeNJvbktL
7zSYw6R9OAQRJwjSmOGAx8bkaOUWckDm0PCSji8qNdBj5sWuRe8ySMWuFGvQmmaj91GNBugSyMhD
DXJxHC0f5gjVUysez6Gt/XzCzYXANUBwDsrXjJGL5nX0j2W2QOWlENWtTKawR0TCC4wcrLGn8gaO
B6lx1s1DXaaKCOZnvXx8lC9x+0iPF4bIPSM8EYyJCGbVcwzXc0TVD/514NUviMhnKgTgGAFG6V97
kObxK/gh9oSZx9AXSuyPlCtiOWaCmvPKglNj+UFc8l9ciPG5yoxQBdRgoZXQtOw+TsuK5yGwYLPl
tqrEeHYis7rK3M7cDGmucMNNLqajFWjCI+FUg3c/HTq1slon70Kru+UAi8Ixy75Wo+7vALuOgcpz
VejIYjkRXWwZNM8wMgMakxvxF+CAbvyq1bIqYsfvKYSfwUWdQkG01p58gR+ELikWrXYEDXiZD1BO
TpaOYOaoWH60v0dgNMk/uVppf9/fpBNrfGn/6EpaV7ZjEQNn9UVBXkc23c9RwOhhbHnq0zzeDaWd
su/PFJiH3tHs0QRFLuUzJae7Nanl7aunCoxw8uAvKnqToTLOOB+oqJ+ohqTpKunIFfQsGfsa2MnB
LKomTQKoln4eD4BRXAmQcNI52hpJwOPP7JiFXCQAY4J4i70L9jyody1q4HdvTrMUztDzpTxCi8Wg
oXq55nT1aY+unyKQCZ1Q++Gpq3VeWTAffy7sAgwY9SVGiA2izwTwlwX5VYdF7FxUoxIhcaiYGqnD
Ouy0F1MxE8XpwPsWCKr6sNvSqZ7otW5as4AFXGlevmIVbF6I0ax6VMQZmZVDw3wroZBFtFKvSozV
cTitSDc5ySQF1EhChFTndyOsVtqeRlA7QNry7FjBKuZqNYDWE+rRXXhvrNgC3ETzEcOIh+5Pzw/V
rPWgZpVtyjiqPl8WRvVLj/7qDwhX4dBZ3c97O+LGMXtnPfSIPAwq0L8VKNz5WXWfOAn1f14ma0HQ
B4SBqX9r5/x3aQu+VdmW0ei26nhgG7QlZrItkjOCv/bnz6GmaWK2Ptxa6Fn1QU0UUcrZeGf/jU8I
STq1LUvsk4occgODddQFT71sKptaesyrDVNuiUDf1DFR7obD9Ni0xmIyEze+tlkjsriucJ4WMYpH
Fm0MXo2bwLBmd1IdSmVpxnZeZxWMuw6DuICmKxdCuoYUTo8Rx1WIR8zVAbd3bQSDx7Hgxev6dWlq
1LSzsf7Ma1fV+E1FvjgFQCrGlph82Ce7nC6NmzyyaMcc35TcqftBKvmFh8gptWdJkw0DO2MNaJ7H
vOUoA3YRCPATvKu2tBBlXgXiQoMy41448OP6/FjzGHDQKS4FVATlo2AdYesgO8y2yyKpz8YcV9V3
/qOHNBGqUnP29D8Kh0OgQYwtL/xPcyIQUewgteyF2Ig0h6/AXOQj3pAmtyz/Wbq5E+9QnjeXR2H2
snxFIAVfLIG0fYgzU/NzSHzZo/XEby5Qw6LydW6pxx0GC6cbwKY1yCnplnRw7gHxZH7+hrs0RwPn
CrV/84/96NkzXVaGtZMiaJKFp0eO3Vo1k+kb865LyCOFsYzw+kL+2S1HI9WsNeJLa8VQV57WuACy
/XBp8q0NT9M7xNRNJRda061/YHPUqm/KlxOWVJHrWne0bli5rkVCRs1A2bGggMUk+QoOvXDos3cX
QRCUywMIuhDwqNCLSEwpeK5BGJvigFS7Duyfih2c4C69xl+9vAL63URM/Ko8q8FvGhO2MxijZ3zU
hM0LyJBaa4IuRuhsdRJhJzcs8019g1ohdloLmGkE43uG0KGOsj4FS2jA5wfaROPwuMIAMzirboeH
u0j+Mk50hkZKJcYNdtshEr6WDf1hM8R2n5pBTwn7shifxSrmvj+O812nE5N1Lzzojpi5VYlKnfDD
oHLzbCM7rpx/2I0zIx1c9kjUHv8jRBGFCWaq6jKBFEJylgXUQsh2jhrz3o/frufBPjlvLyHNfIZq
kmVfSLEORh+hLuiHD6vvlfjmNN8AGZNbr1BsAxrGGGVIMgqadvwRPfQ+2r5sCOckY0LPMUs4jqKe
TZktS6m8MA0XTSRRY4/mtb/jIq5Bg6RldkwEUWyXi1M85EVwTxX7907lLdV1WHkN5kt1RjeMau29
1dMF23fe6/BR9/kixg4P7M8ac6wLUflDf6deeq2E+o5VqL908lijlsYTeQOlrp9GbTJujs7f2xlF
triq5EZYMtOsOlEJDR3hG/Gw8rjHn8RM2HWz9jbqNqx8cEW09uP525JX0qy8Psx1PuDOkNEg0Ebv
i0E5U1TW+MGU7PwB4cvG6jQwGQ1WnTo/59EKwAxhJ/6fl1Go5JyKWD0NXR159Wm4rboCFd3Gx0D+
VwVBq6mT2bXtHi1v2JSefUsXNZ15C66PHIZUl8iakqATKwYBdCmlKlJEsr38gF52WCcbNDLx0l+/
LFe7Z6BeVYaYPbPVYyaAvCQ/dZ9tUZLML6QEyVLDYC8Jg6EpUyb0jO7RuZQbnAe/PeV3afR87aCI
F5GxrhmadjmvY3vSoizciXshnrWDnRJAZrCz69pZ7uGvE1g2l/CF2rXNQ9jqjoytNav6CNIuENoL
ltCe8/BzcRCLETCiN3gWW9HBkTic8iMeVFBPB5wJGH3SowHzfN2YqcDBcWx16uquHgQ0ns9qnZzT
vIxIseFGyza4anm1bEwawDtLC6bSaGGZO5r9lMbPBoLwSZOnDwIhxeyrxFX6C6a3ws0foWA79bGA
UtyYzYQ1euyGSMatO8T9gupx4vUrFfZgYqW6fnwutNwCsazc8deE6b58kDVBxc/4M85Koo7pAE1w
8CvqL3aD+roIlYtUHZw0CcE1ACbo4I/5YoZ5PtbhDeQYyhFKHkm3R4jbxE9zMM/528PiWEezVqdk
5zrtf9jspbjIJRnxva/7r42tdaYcDJXCnjtd+4js5hUvF3eWj1Rb07+HD6GLZ3XTsHviOQuMPMnu
rw8576vpKrSb/ijPvouRqJNfLzwvVh/OnAaduis+/+rgBTHqgjcmwfseHb63IS/w3y41Mrvjyei4
AuXkUtOnOnlfsIM/gxovm56I0bR4wYOhytc/Dh55LVLl456Zu0BHgAid8PFQfZ5cG7x0XxzNcCme
ZNsxU+50rGkoi7+6WGz4axh1oulogWqW6x5KZU0B99MQoWP4VW+Ryk61EE/1f5VNND70ZgnY/SPK
mpYqPjZDUdpTpVjW5Pij2verMHWfGoeRgy43oc5YbQzqRWSYQ4kWsze2aKgJFTbzjiPLkFJ1bK3D
oco7u+dTScMklwK9j5GOCsDFX+6BvhbVD3fI1vhmvW/wLmZkOAoEdpE7sv4DVI3/z6QDxPcL7N4C
IHhOwnYsxBv3eyEBHpHyM2AMb8fd07pmwPEwpG8su4HiYgMF+xFSDOYt3zYq42GrWTa8zDmhDhlQ
g7fRH3lPcSmX6XRWdPXm+JDmsc3a/NF6CR2HvEFMNauMe6BjXCBfDThtEvcPf0H1bcdosr3qLyvm
dMH8VKPJD1KvL3c9muYp+LtZP241xW1G/OeYscTVJyG0/nbydRhVakTZJnL+pFYaozSjnblj9mjB
UH1TAq6h/WTkyQGUbkIpdLJgPzaWR7anvKDUkRq6MvNL/mSx2OD9Es7q8REFKrcdisRkQgCN1jvc
rk4HFbCb1Ud+zjLdPl8Tei+zCefTaegQX/DhLD7o9Jpl51HTXIamW1mlG+nelKDvXRYzLlVfo5ha
6Mb+gABdd34zI6SyqWB/WSSquhVjoJmD4ZUHZHeOhx/b3z09S9iwCyeKSI41S3W0IAQmAjHZDi9a
GroqUP/Mjs+2i/YZeO85uTA7WW6x65AdinTjakaVOACMyHAYHM6cKUkRPbraZs6h02T0O6t6Fuyt
4m0DM5s5aLDTEVu+mjAGoOg6InHcaOOrqOJTnIU+qauN+GG3EVLBWl25RVdkhxpXjiGCoRS0N/Y9
aiOjw8FDTl15WslRrpopyj1tBVje3dL2Zb3afpC8o1c+oDXdbJNbBl4l5Ho1/xQRVC/im/FdkF94
O8Rs/5OgCqOamKZjW0eMsjJ1viBzkjA2+ZPHDhieIiMTdsDVqikbzPd4EO//TphyTbrFhZ/egQcG
UG1da/++CcO0wGd/jzNrZsSJdvU68rKsV9C1Ycrk8H6yM0u8giRUvKNtTI8rSGAYySw7PqKJBf3K
Zym2WJ5CqPWjPGVzdP3Byt9o8emZnctvSFWcRc09uzGHEaWOu6dMvl1mz2LAcL6WxrzGkolqr07W
Lh9H7x0N8d4SH9gXVeXyAK1hKamaREblTWHNrFWOoRUMwybqWN1yg6civkh5XSZUWDS+SDc+hCuH
mbuJ7DOhOGUcl39cILaI1Q+rjyVIBenTIM5ekv1PgF0BgohZuVcCZkn46jYDcAfHowiQVz9wn6XB
s+xVOApUkNMhkCTOpj3+8AK9tQHF5BZp4R7u8Xz7kJgvQL57ystjuKNDDVPKxAcJ4OkyFfLkrWzH
+2gU7Nr21VJNK6UmermfxoV6eIBTyZ1m5xw2ysDt0/B1+8BDLNJ73VMM92E3pE1nuR7Oo3NvVwuE
VFH41UKPtFvH09ZCMPEj3swd3LglyGJGEPZF+NQECPR5yRbRGn1bpq0iyGhShdVz4Y+bNeyvhJhq
/NZe2Urf6f000Zi5KdBaoanzpI8j9cebPcMGAD62SWSBUfiwtfeoXDp8FsCLVD/ne6PVz01AmvCw
y3pUHXzP6wPXrBagYFn0DNyI/hV+p3keBRWOJR6w9eAOFFe724CiEYBymalxHs8ePE8zb7zNBoWr
hDIhFBz1zNY+t79TXJwvsRjz469JJrV2MBAlRqufMAVdseOmQlgphxY6VhKpSkjCZrRfUmeHSrKQ
J3zLIjCyFkk4lszCwrG4ZZZRA4lE1r8XcKUy5btWMHZWBACjpQpx1DgNNVkFtfmlaz5DL0GsYdNW
ZDujXfMxdJgzbGyYUev8d9Nr/FLZajW+GY+skPDJVKgvdMovXWpgvoLRcWeENybeYLVjwfS5Pw8t
0rgJcVK3Roy084eohQIw76kf0p4uLfzuKfJ5SBnm7OZqIDih1wvqB5IBiEfztGZKqO7yBm/IC0RZ
x3PLkOm0CCaNpbpU5KX8NnUNzdgv0VvQymBYusKOgLWvuMHfNho64lrLwQVQH4ba1z8l86lGwjqt
k96IcEEgxLD1RaBglJa8OGACrKqtNcElfsWdMJ80ANvZbsXBKidPqiKFjTparHU/ebEyIMhRVYul
BZDZSOz6hp/MQMztltG7xUTaT3jHnuGxw1MK1DCgtBzIEAM81jkSiB7QlmjKv5nn+UXJ3a2Oeqlo
/Ahj4TuJg8FOT1r/EkpMaPwfXE+bvJO0O1ZmIzg+pA1ZFAbNikXu28i9OXexgtOXWJ5sIeMSY6br
HE0Rz1rm5HNIZKpfiwOhf4yXqGUhNKxt+58a3j0w7J0or91RwTc7S8VetSikWrYyg1r/xbr+bO4p
aGhOxtNOvHL6tiEyoiti9scZWxsgCxHdALo43LXE32EOMJ5Ie0Kp5EowPCIVMlM6wu9toc8gJBWJ
3Wc5LGlLBSaXdaFVmd4doERPfWNkZ7kUgGPQDq+lXg1+uaEm22ZC4KFKxkCxmEXHouMuY+zrfTb/
BRHEKE6HejhLX8fx+3GWMCwYhJDUeqOT3W+ZgnHZfo+tPV02Iku1sF1diwW5xEuPkQmVvc9XERZP
IX70gNeThwcvZcRbOdtbz7TxMamQzAOzzJNH08+dz2QVmyxVMJaSVpllXMFDHl/t+KHwfCoqiC6j
HvWAzSB74LkHxGWnHZk2OA7JelrHWZ+CWWAyM86MdcGChAsm4stv06ez8wvB4zEkKcpKSRkJJKuB
Ry08IK/2mKCP6WKxq4VDQrxjjPxiAFenUzTRkeuAIFSXZwrZwxzByED9A4aNcgtxfmyFjrzbawfl
MCpPbwnbsBJsOOMX6PX1uNFkqF2x2Zqw6wtNAefdq/QSfn3yhI8raQSitou7PhuWKhWCxKhUaWOB
IgV++UcK4+AOQcRLrLh1ahw5oDZlPBtqQIebfbN1bL8Y1qHAl8IsV41FbFnoxSbPpcRwhb6oYL5G
U07SPDs9/JxFUr/0YEEG35fzbRVQu8BQXpBibQeFoLq4Uj4HhqH9ukR/IMheR63n3rqfExxH8iDS
r5smXBigUkiAUfIYP0/Vh6aXSmL3ya+oSolwTGmHa2PVSJcn4Ug8h6CvxLNfYhGINDYfl7/n00O5
qnesA7keeb2gBmjFeGhV0rsTbh/xVWS18N+rAEY0649AfuTIhv/HYlzBu8qXYzLUjfh12NNx1vg0
vqe/5ZTgxIjSWTX6gxzsHMvQranV1TDsRZN7/C8pUCG8spbAF2ljt73BQa8ftut+rrYVmlHKSbn2
l5ZcN0ugQzTHtG3+FRBy1ujStsvP9XV6bA8EOf3UTlfMN31lblTKW+LRAHXydb3+3lsRaNmvDbxo
784OGlNKj7uuMxc1EFkoWHTuPeOfSojONhaUd1d+P38FhPSZ8EZ88/h899saFvdimp0F+eCaxuPc
OaMt9MwaDW26RcDxuB337gaXl2FGYknB7TpykkPFAwXXxrEr/1KmLnjpCWpp4VmAC7cdANjAU5DE
EA19pFUuB2CZX1BXATnQ5sFQW824V/M7cjFGkzRxVkVsoN+NJo6jD4PhhDmgtXaOPY5V0ynjmPkU
4rjyIWfoOFRIgtLZNF8DFBbeWbT7lpwkop+DYan129GkFqXa7bAzncg697Qm3jvx66+fyZepTvQ0
yesMlmj+XrWh6/rjTeBY4qah7l3ftLCCKkg0aVS/f8q2/GjtCY9LgUiOQClCvkVJWBVW++SMRU+x
Wr0ZRMIGgu2RSH+wY48qvjlGzsgcNPhPwWPos7iz5aSi9aull7QGMGH7qy7m1NN5mBrByJorVGd5
4PHEO8ua6pNENUkzDdhUI3bQSsENbqbGXwgiNFWxNnMWEPszLNT4Q8yf4G/l+3hW3L2l13X37AuJ
/8s8SWA9yHJ5edb+gxGVIM5V2KM4pvsyYRsSgro3dVbUMH1ELoolMcFTxC1DQsAYGwtFqswrjXPX
5hMEQUOzTpiSQOZ39jOLE7GmAyyDpVsFklGcJ/391K7k/1yU7RBSWC0iPKnJJ5+T/vKBHDJYsTpI
4DdtPmfwNX8FhGDbLf8lTC68JySBCsWynHTAw8lEfsIpuAtBaMTbLrmtR2ZyaOMPejkyww8Cs0Wa
jAPLqXuDt9xCeGCR6E0bVfJ7iiUqIUjevjgRye1kGfm6WGQg/LXJ8jPZvZFj+0oKtc6Ikw55MKM0
DA89q9UrFUxgWNgQuYHkMPbYiYj029z9vfydBA4RpRUSaWGWh0b6zbnXyEtVPJIGqWFpnbj+sEtA
qrauiHYuTWJR7Wx+KnRNci44ZtuDPfvpdANFW1P7uXG9/PKPNnGsPzxuxmLxhzp+ZagEmVsZRuEa
vVE0l/cJPs4F4QHgvT3WXmj68F4NMTn9PygfA+O/4XP36QzrOCnqIFDWvZ8Pm9+SyFyMhOH2N+Dl
Be2KplA7DFo8Gr91NiiHBqAkoO1O322ziKTiOUrHt47PvghGAiqC34hh/AMvg+03fiB9sVbf/vC9
9umMg7BZFY8R46zDcQr6kqxjvor8oIwgGLMQF5Bb1bXl7DMMKFB5ahES5/d73AOc56tgFp6kNITP
ANH4BHUDBk8xvtUGNQckeju5YkNXFhnLXVn4yCZcUSRBJugm/9wzVEGrRpj3yIaIB1ZzkwVHjIqZ
+Yz66hvA+sxjdG0waxAOBbA8kQ+pSLpAvkTIvFk2c1vk/pUBSXSl4HLw9sXJwoMk1xu60ydK4GMp
OW7PRbiN+fYl49dAyYu5kPn3uC7CSFMcwaUwpm8bQtCetZWrp3Wajr92qGUlKl+sW5o7vcSrAswX
iLJqiaF/LtZtZerrgOvspu0kQXgVKgmu0EIbgh/qGUX16c5cmpwDLRbwmyYPpKt3d+B1/17FSzX1
P5JCbGMpupKSfoMMN4wEi6Cww+GU187j7JhVvhkHRIkDPkpNV+kWq4J9swgHPLNpBXZLtL+iCNd3
5S8Aoxvx694hoFZjW4mhpmOGEef0VsQiBu5UubHiXU8fs/XjXTtWAEcN26DETjHPnPYKcz8frc2m
5Dg5FuzThgXuLpmQSt+d7rh/ngabfMZBdauK6/hN/gvtvoHjS0Q/fzxDZJeyYhAuBEAQCWzuAV1I
Lzo17qRC2NrP5oA9ksLO/NgeizWE+5pbmJXE74JTv1fbIvC8U2KJpQ/NEmgLPBhclEk3LmYVZp8F
2/RNFpGqiaQt43OT4Tv0uIEkSh69jH4G2h744iOhHT2U+ODfNmh23id8fHZq5ZrgHT97mhmEzO0w
KfazhajpEwuIuKlYs99nyVHspuMyARo3u4GnyiK+K8dkgLG2OXXsoCa0rqOIOFibDtseiK6ZzE2n
UWZ0CsKKpWpWZnfY3U5m0dNwfu+BzyMnwPndaZDARsuNXsQ7o+dfVQDs8RAsT2y0RPm5qCzv91T4
Mx3W3ljdqW1HtusTB+jnDBXvNTt+DvlPMOEAyv3gaNajJu2O8aKW1pRse4q8tqr3t/8ey59IEan3
fLWAFo1k97fUEBdn+7MvCRBhtr+KfpGei2hQtBJiH/SfeS/y3GSrMCnhWS6+DrHiEQ3AC+7sR+Fd
+ZMc6PlUaEgpoZRCJw5WujigdY8DPWDMk2flQvLXdKPVx++6vJuzlwf3b7HWVLSzb3jRDRIpCpzw
2wn/t8GKkaRJeuaQc22X7HsHl4P5soTTNNIHOLZfaNb/STS24Qh0oH+kikjQ8pWElde33AGcEDjH
guzjfSSl5zHLohFTM5Um0jgOOQUkhvP5a7UnWPtRZgvJG/KAE9oifgo3s4UQ+wW2e5+iRsAHFeDF
k9QAUmC1yYO35nVdU+FgowyUzKKo/diZdrm1S0Lt9WBv3lPRqI97HfnacO3yC+WtYb6rYpO3gkfd
VLx23zX17bzNq2kSMxEhOEvJL5dtGKXWSfgNrj8Oqbz8TfMTqRJ/k190TIWzkcBSLY1ITPllfcAk
5oD3sPZaKvLwaMF+MtcGZ0rrVUVhJttC0KnpnSu0BYZbhNMop+U25SXoqFI0Gk5R+/me3QDVW9DC
jRB153jYix6dqa2/ZKFE9tnw75pBoHCWFy5lDh1BlOWRERx3mRFx/6sISk1qO1JgjdL91DZZSw4R
GU1s5VsswYnEZtZjno21xwrfC3Ay526jWYugRg9N7D2k5hyU9mb1JbnsLBy4LlWpq2WXaol7tM84
17eKFU7L/dAHl7fYfkJoL5DhOx9ioDRUH1Ax1BAg0EDNyrwb7RZCOSpZ8ZO6sxq1hzUfsnfTzzeY
NwabZxLRCQh8LhLbXnlPmR5kvR6fVAjPn5iOx0TIuP1PR1mvGIodgbGWjhmyjHOl3rVlYKquN3dY
XfN3PAautoBWJ+Bxhzp+mGclLEPSbkHG2QVIEWvGOvwt5bX0tlKlahP7z6OXT96mC92degznNdMA
BgtsQofMs3Lp67+wlo8lExL4m8RWVSc8rtTUR1TnF6chSEJhyrsANxJUANDvQr3cNHfoc/aXOUDy
ESr9CyNmo4IGzX3jGwlFcLN+6yk5z7PIvskR2ebhCmeZK/ElQ1NuDHQAZrY8Tn8IfueuYLMuQ7wr
Lrt3b1qhOgYc5bFPB1tnlqd9RUXRWdDW6/6PfkfdfP4hE3Ug5TJBl559AXMHDDkouZPmOIffwTP7
x7bJgWqV5iWrXBH1nspwlVIy3E9mplw1n+ONZNuixBu7u5JBXO9FIj0nIEji2PEPvqYYZ/9ErxKQ
HrtDUBglm8YEwL4hMo1sI99hRQKZ/h03Rk0uQwXwh48K/DVyH/RCILAz5ept/skDJrWT2enBiTVo
zajgqQREv8vkM8pU5omQsOVwM9iyNvgbW2PhTSAUDMYM5UVfnmPe9nH7nuNdRbH1nEYwryshsIdD
L7sBPCguG5TB5IfLoIStJkDkgAiY1SfrDQH8G4k3d5Gb+ngrf56OjLZTqxstOVbHN1WDRbuCkl1D
eiUMutd4nzSCi2OPxZx3qbYN2I9p/JsXDxMxm7tuuYM6u9FSjJ1GVy1zxSUrl/aHVNV0LA47Uxl1
9FZHo0mILQ5YwVXnzWVOyhjASLHUUTUT5/LZycQBBgB3OQ5419XN20lEDN3JdJ4WIU/W7ugGsu+j
p7J4wiQ+HGQrA+LZLcqRxiqjWlbAHOsYoWpP/gA9MDm6sWNtQEzNC4pILvqGICD7/LgYeAaduee7
uDQ/DDW6BYvZ7fm9KG03IPNlNWldZ8f4cyOFQIjq4WA2kMwTv7GdDC2URC+mWycBLIczWjTYRNdp
ewbt7PM1NQSpuQt2vQk/4ACJB2bYtCWhbr1RJla8MaEUzJ9FoHrWmhswURfIFMtcbG17K4V2OIlc
OmLinTPwgyPf7Q3IEMRt0Kcb3+ebPQTL/Y6cFEherOAEgmrak8gqph70u3YU+qz1bK0C4iH3AHC8
KsYob9LGCMbGJPXBLKU3uB9mPEi/Y6f24lkGr6pGjKCdZO0xWKyTRQV6tGHiX9L//uJ/ALWy2gdc
o4qmH5EMdKB1BfpGhePbxi4LY3rmGBPJURtIpbFPYciP27q7Ez8Dz9oTWPTMDR1e2zoMgKe4iWhV
CgECDLDn/3MneFmeFaupu2qFfpbQwEoZT5G62HuergeZvkXYMAoxOhGpOe2zJUDoQg1AQGjPg6AJ
qEmGA8IciqcwqWj3nKv2+PRUYURW8jfs2SUiLE+ZlgfJ1Ckyc7CAtIxJKcHrJ46MsVssBYM600Iq
70PSdqeF31of+JwEngvEA3aahTWVSix6TZhKma8lSNoXp26xbLpun5dYc8OJN+wAlBg8AL0NhwUW
kICOKBFtVqf+t8X/kAzG/m6EF8oBafwEghf2lV6GjSMo8NgTTOTIRo6OlDZPSJ+KQuC3wYxxcq2T
sF8qFMOfvZuEGFwmmpKZyA0JfTzbwasBR3dV/ccMA4jooirylnqAVncBzlXJKBuDaL65fM/jgIPn
PLucHJHDrE5TwwGsg9Kw7L7ErAIGsibG0HAVktr7LCmaySvzVDZgFrH9w8GstcNP0cXx8u7mzP87
LtqTpkRrLmVhCPr08TD+xlBYZ5leJSNc1CZkBIWRbYnpl5dU5s2K6ez9cJwW7bYiCOaP0/G+4GI2
9xz9XQohLonqdy+fArl3Kkk4Ob1Wvw/ngp4sg8vKVwJDufJk0LY00FW9SKzLSbZNEr+vgcKQcNrI
yejMzw28IliCOP3xwb86Qbn7D3GOzgKngcp3HdMQFQMqxD19A9CZcTbqhlBSCIno4w/ZuKMLbWRF
WMoxnvHd59c5jrkiKXXtopiZe2QNCYir7FWfh64PhSzgi1zWm4D6Jko0YaFn5tZBkAYhohvgpaq6
E24x21lX7N36pYVkEEx3vIEK4lqXwCKqBfu1lSnCxwxDkdKDoACM+bF/uM+lt3B3MG1oIUnIjpRE
+zJdnYqEOUOsegacOA9jLxb4RaJIOKHlQWFFvB84e0PQXjbVHB1wYdLOEiMbnBaU/bKgLelnCcAv
n9XmbFhfoBTnjuF1WhSRy8LmxRbAm30IN/s73tw0Cr22ZYRG0OKoRHfKNKQKCqM0DTBoF8TQGVCP
5Sk0zxdyHp67TGTx8LHgaOodZr2s5meiwZwP1k4HcovJZW0CQfmeq0ddDIZkXy1lSVjRapE4dggo
HeKQbtrm/3+M6nXaxDTS3JgT86rXWgWPeK2kQUUTum4RifCyDGchTVMSRZSfJRqSAaYuhzi4ErhC
dDPd/aWfCwEw8K1PA/uq8luthvt0TGKfiN5FOHkzw2oOXWqYJWo4BXz/3RTqSl2jkkR5eVuvfqHA
IBNzX6sxv9conJqiaYMgzEl9RiORkSB8ME628KVUKv6yvcWYSNC8J2eZppT3R7fd5ALamwh4UM+H
sRC2RNrc/E97fmsV32dw+qLI5FGA41U1elSH93iZNubjt/Ts4oHV6p+/5CBhq4VEcGyS1izJhYtt
uQ1VGjTWNzlUrlOkrZSOKTe7StEj7XBGDWuHd8ciVc849JCXcbLH4qB3UFNFEHIJMMDA9Dlf/8RO
S+ryCLuWGFnDLvz+HS6gewjtkLVEiGziEkr4hgV+NHKlttVJ3z/X92jpnFupFoHsfAjGIVkWQnU2
+ISOo2TrhsUZYZWEcWIrQCS7f5DmZxTIX5NDcfmpZKfE6AFgznTueT1ZldowgFGy8J3vvhxAvHIA
NRdgodIpcpgc7ocNZdxqUZG64G2ePfanp+XS6tC4drbhrpzeJxQKi7D8R4km/VG+Ka/sctlKDl8F
CCp9V9HZcXuBsdLXLRlRihzGRaJHw//7/5Q7ookt+zz9dWymAJmqMl3o03yzAfUiE9lL/ktIZj1e
6WVoejtJaJHpsUvgvBobqMC9ylmbGFZTMlfYIaOH+jsog4wCYdwiqBUuqYG4dRO6xBaTT7YURA59
+DVPvrAvK6qn7Tr8BL4YrEdlCD79Dp1MjHXS2v0Kni7+zjpMuqfPQ9ucb7XxKTTFPlrRuf41rYpp
L4hoX1aPn7iLBN9uOmhFSeFWiVeEgLi474FzbywN2F8fcq9YO2y0aP4d3qdEk4euwo2KxwRTBB+T
sikNrdkp4guJ10m1cIvtwMWQYZiDeidumf6GHXz/Mj3ZxHx5ytCzWbVKhRqS6o5e2P6xM7R/7iAJ
aY7xu8omyZ3YFU8Z4yqMlex5taDgD5JD9uRJUbMphwVhd66EbSoMb9Gj+UxQc5Bn7TX6SKSSyxo0
+z4FaURtsOriSKgfndi+s0XJz3AOuXzxme7C6QzSFLXUryJP6CfEAsuTbF1vNVCi/cjPMb7zSSGM
1TpVyGmjH7WxkZlTnS2dYhP2eDbinS22x1Wdu/X2ctdmn/o+XtzTvJIYm8kfXKI9e1w4NPfyyxX5
NxJhtWlAU99g28XYmvkYT39QGANjmlA1QPufLfIhcpiS7bIoqTi/WG1h2NNphyg7RGuyH5iPxNMG
FwL8OIx2sjUOum9e+8QF0lmKcAVf+qxogQLdoR/TFPbgLf00kWBEAxvu0d+owM9XNuJzhic6BmiE
HfOyrZj7RObVqtvtVoHkkY+61rZvy98jw41xZZxbY1Y8F8PF4EHb63ASFzxlYn0B9END3wRj3/Xz
QO1c24jeEmCb17bp/sGZX1mWzxenjcoqQ92dGrFaWXdwhf9i0WBfH4Hl8CRYCM4Diz8G7+lpgC3T
rRVFLnBcfjxnKSmh9/a7+rZ2+S9TCzxgGGCFrA5QwPEVXjaSgkQt3q7Ew4zz1gDdGnZpqgZR8dLF
D5qXkRi71MCv4i5YUGeGyQPwXmkLFxARFL4nnPpT/9+0TIW8LEant7qGQzFS0ueWp78mT7Db3BvA
Ehi5U8mmWYIlBTPzC3yrJ8SZXMOuBhE2nUk08ka5l9FzEvH4Kg2IQGTL4FAoIzYAu2UGJ9YY20Cl
/NFUSc8pORRd+CTQjTGS1GJTC1oldNFJOZjdAz4Dq9/DsLd5ygTNLegFJd2f+Q5QngAX4atKESeo
E3vNxVYHp50c/f27XiJ4q5O2E++/vAY+r4zolBATRjQDHEtHwLXh0ST6VpPH09ZTKrN3r+6KYO5t
1MzJifkgGmCsfR+0lVaSoXYZnxuNfiOJj3R/U0QCOwoEgCeWRWT9LNw1WUEAuQCE5oVAC6uV8irR
lEh1sLDuIAimfClKea6djWGilg76viuE8UlnlDiT2J9dhAj7KxGigz21a98ctJscRoS74FnyC0sW
F60MIQmiIhDnwcddE5NOHXA512iVpO5njA7OJZS2ohqZ2gyW00rcEJRaJMTYE59883kDiwrrxSqI
roec1lZAseOOXsu0LoWsRaEz0paeA/IzlIQUEZYne5dw0d0lALZ4CfRCYSmxMggMJFXf+YrvFboA
qQ7qio7ITOdSZjJsXNRiEzOCh0VSfZgHlNRmoAgcihdeT825Set0X9cI3nOJdOO8crhvkIGYk3TE
jVTuKwoziNBOSQWbwXHZanbsieZgC5viN5VbFzvDh8zEA6Z7bap2qrwP4C0AvXgivCGqUG7YEwP8
SFcOzqHr+au9DzfK7qA4jBV9Bx5tOWrZD8Xdf4DzLQelo187DHaeoBr9dvXgGu6Gmk0TvHrTS3uH
Lddp5diL8FzDsjbW7osCX+6j8uRd3MLVv3eChgQxPnGwJ2l0kLH46BIq6M3Op+peVMX6tyIfA0hj
q2qUMLlA5h2Ir+YiHrtc+Uzmsxf1evDaPBKV8LtF2mQIw7+Y5SonpjVpfLJUrL3/v/Q/lgUfIFZp
tjvyXJvn1Mdyff1m/suEY7w2igJQhPyrLZ6o75gIBP1YVWQx14ij9lBfpEjLN51MdbT9h+cSsBdq
VhRlMQ2ZNrMaTplLuGiNT/vUOuw6lprzxMaIrN8mn2sPNrRobjQRMjQRLgmqebS5Fp1B3qHWBpsw
Ojjgra7EJd4Hxpylbo2sc8X62Hc2hUFz682W2RgekWDoW1mUPp62Ww9yez3/5uRq0Xp2lfBHV7D5
0tWEpEhl3BfI2sIlYXLp8JQ9iH4gP2UEncBAOFfHfmPyVrP1oKR939mcmO0d8yhLGvaf73LI53Mt
ibrXdu8RANaSCEuLjaqM8eXbmuGE004OjMEYA8M+OExt58TjL/iiusFDOAdP/k8nKLxkFFo6AJI8
8oTE/EZHDFRZU155vxo+77yPAr2U/G4ws//bX2ru8deoiuBBeY0TaRIS+Fm4D/B7wjAquByrmlQf
9KgQ+zZgo07Ciunv7Ld6glYhTx4rVWHcbUYzw1Lf1bL1GNGqcS81Awra03HNmd92MYgRpvxBDCVI
wozf8yrSEJSatM3LX/FENhtzwg0wPGcDPsNLc0CtQmmTgARvf67URVV18J/DTAiAv/PHF1pM15V0
O/0xRGXJSTmZryf9F5oqdeb5CuKHKxWB+YK5miK62vX2NECwnsCN2EqutsS8D/PsN9m96u035Uvn
Cwki8QLDSXjXA/7//iJijM990PmTUr18IejPOu1jkAFdKJX+c5ZvJaA3bD2aqxWD1XNPdy+T2/FU
gcxhauund2hED0rcZuKv39mYANmNsfe6e5DKIK5Amnkf7uWMlR6bmN7Xz9uP3Nj5IL5cneVnqH5U
oQkAT1tGhSNolLBsiVEjTcXc5H1HTJ0st+IlxORolwgee1l5OHhzh6thUJ1DL3itFIp0OpZTiXLU
CMyX8qiCGwB2WkxqiLorC/7kRC7v/pBTjvcMr8rlvIqgIV4KLm/msqPLf9NZeNuZeoi0V5BnGX1S
Ln0vm7YROe2lic4LteG/2f9WVzYKx4UlsJ40VDz9t5FoxMpaBF6nZDJOGC9/83CslpkHVM5eSUJO
R6qYK19PTXH0IPwi3x2iosHFOT4hPu1XXOwoDFtcsK0wa+OPcb++CbwTGz1jAnI53/ZlCZEtnyiD
MnLETCx6iwaIblg7F+UgI5VrJf6yQCFMhRIBNcbZDjSBg0zSdx7/kMBg878ZJNJkVp7EOFBF5a/w
lmE7j0RGyN/mX6t+S1kGabvHW/82LvDmpPT1vprRmRHcKwjOkS3pTFMZ/Xae4SZ8CiEeuLDK4e8H
NF+q9O2jdNGs4d6PWMYTNQNNEudqRtDwetY4N7JG5ete1zXaASJC5LxuBgr+EFE2qpzdSvIGMsY/
VmhDKHZq8qjgt2cl33fvZFWEe0rd3cEMHa8BmWE0845I6IGqvpGlK/1fsvdvVnm/jYe4azLwVkzS
yBGgT2YLZMy0WdrnGFX0+vuxWxe2qo7uHghu3ABMndONERIyLKAM7JGzDKaK+hWno/salkSNQcO5
2yMoi7+KqCuOjffpUkugOrDhhWZnEQyQkoAXXOgPPJkdfhCg7Ke1/ZpQEJAPt1B6KcQhE2O+YNFp
i3HMR4FTJqiW+rpuYAXI5ToAIxdqwoflPmWtLOx3oV2ML2SqP6ZpjzSxkwQLZfrZvs2EAmhlt8jt
tYsXWoel/bDIR9IDsSJh3royrSIXQlfhSqwLyo1hK+0CtFCNRlnsSbkF9e2lSDG0XP0nKgSY0J43
EqxK/vXB/oS8ORsJN3rTOvcIrTmOf2rh/bAQ9ObKhNIidTzlaqo40uAnNt2XcVFC92q5IYiK12Rv
ONnWHBZcvN04o/JqNkfqEiePGUgSNxQroP3YupC8+IZxEck/ve1TPP8s8GZx1n8Fk5KcemqSXI6l
4IUptFw9PFAErT0vLCqZtt4tV77xgDsNnxg0ogWEWTpQC7kVYSgYGFmCZNiSkaGqioXQmQgNEn+S
uDkBZ2LVr95ed6lecFmRkA9qq9UaDw16aPf8sWpEl3xenVCDeJ22lqv8ZZs54JGMP6pgR0bqfUt0
B6PBF3r43XXu0FzZXHbSBVxNsNDuCVBcQtjD0dISKtrfHEjit3qtjXe2fYzAhMLdsPStbHQPi+wW
AdD+lNn8LrrE62kPz5El9xUMoPBts4anXTGFEu1A6GhjQkO1JUPzM8zw1PQbK9TWi8ibI+2g51e1
MMm6L9TIDVZliGIjsbTxu9rj+Q10ncaKqbY+dXV/9vLgy5xmZ6pXvj9PkKW9Ui9RjiCCXjV3plMZ
uNyEw1qMQCtg84HCpKsmvGHgw68HdwWFQIL9YSCsMtJpH+i9ZHAsnb47mZQsBnY5qeHg0t/MorWJ
3gXheKaoY9orBLAiXvMs4rbb1ghDDer3Z66qledfcKwuov2KtIDsbUvip4/FdNpZU2gs1qOVPCQC
/JNMFKfJgWc//flTaJHv1ste2/ctlgUmkM1g5xzhIdmNGQ4GCg92e7TV/bbkP86q9RP85G4oLKbt
SnJkRMz3P9IU3VrbWpdp4bEozXSirLJ6zlkAzpwjsuGSkPz7RBi5P5fN5dqaQY6lebz04nLMY0+t
bgFPKaPBfV+oK8Sq+8egpodpVbu7NTd1MclnN6YS2ddyEPTB9z2cshyInw2/vA8+HshbpOvMa1Yy
3KS3IA9zl7OUracrsCzxKxT55rHNZ4EmkoKE2zjQlGnbzXzACIHCtDjP/gevKmnwxYNfSOWX5hXN
t4N7kf6NhMC9+WnJzzlH9OfFtuIOV+ixtvO2e6wCpc6ge3ScCmzUTzA4rtQ+eKURG4K7fAUD4QON
Ro2dAYTV7cOFI1SczIkXP1l1ujNmXkOw3XB1h0ERkUYpg6SfdFXSPtguAkqyymX17kThWnF8ev4k
S2LNeeEhtfMbunPc+zG9e/84vSES+mVbEd7/jpzyKnb7wkVOjQYVLDNsETyJEfvQE9f91dSZcFVW
rgKRO9RBuVUkmgMIRXBrVmo7Esq/vKUq6s6mVxs9JRp4o89MAqdibhCOE4BtZJfqen5w4QuFELPP
zT2/9o+vRumM83pBl4NEzC6xb8YCY/Y1VAB44BF2Zyy8LQpKhDEYVofHTeEB6wzcm+EQ8+TtEneL
Vdg9MJxfYqYDJaLlZeK5chQELlQm/+FWUD02Rtz74idxE8+913f1L/SSKfUTrEL+lj38XzmlA8q+
oUSaGRMwtPqW2r6erfFS9tcmxoYHbWUADIcz+BWJNrP4RVUwTESm9kvjUlaDPb1QTWoij/qVsrju
3C7fqNTb1LpkQfzvA+8/ciDHDRN7l3mMw113N0XYWSoH43aeY1kNmZdcDYXzV+8SfcHy7seT0gLD
YM0ckEa0p4iuSaUvJ4Y+Kzrv7duDceYBzkflhhOCfUXh2Z48VXlZCgLf7AoRxSwvlHHSw4guJUKu
ckjWWTw+xcXXOvK8ABoHW0LUMMiIh+l5lVWmZTQlklaF4fdZmBGRd5+pWG8SBVH6bDop1mkk2RZo
y/UpmoxHEAzd+iY+CGZsVCVBsfKpLNauPwPtbhqytHoipoDaaDpEJ4uWvpPq3u2ScaKqUnE9aJcj
3BnMn+BG7cgyufczXOD+5+BlNOcUG+HNjncnkDz/0eB646SDZUyoYCWyKgpcQCDrgB44IR3jkb43
YLwjhGocAr7Eo1sJPRipf12r8UEGDT75qTShKfckv/BmzNToyHH7iMW95lXbbF7lBEZ7sClqfnV4
DKowrwm6tG0jPxnC21K2m5POeQyrj6KB56q0Oxbol7NzjEaNbnxHxMYQBfCfzkIc2WKy38/ezYtG
twI7xpjZPq7sBA7c1Y+5LS5vadF3IUjx4SeBra1FqkcgSRB3omIrNTGEFKe8lIMbgjRyG3BOjw7f
f97jUdjgKwK0WvSmWhqRaoSEmhMUQFH8EJl3vkCpANe/9KCJybnNg8wBxgUXYDHFY6XbE2hXUvA9
3HEs+huUtWDXnjOCwOhnvka+/mG1gU/TYaBmnC1B9yECVJFTcNyoyljpkFavRWvTWWhj1NvcJG7K
QvdW6i7wPycajsF7rlCHo4+mbMfVZO4N/TRn3xx7DFhYtNMvjZifiMb7v6230us2ORosaB2xnPIC
RG5tstKcf+nEoRfSp3n6o46FSLFp8dw34whCqMTO6HKULhMQsPchh3fA3turJE1tYJpvBz8y9fs/
mXMM5h/C1zNNMwuwWC32vpmIYvdKjccqx5F9/X9zYgGIYwwJBDvE6n9ikf7EqWLfbo71ca0oxXrY
J+9C5rsvZKU7WovD1AMoS7Fg0zBnTVnXJBxWrpjpSRScfpBKVTcpnQ2339qACMNWSEdn/z6zCPVq
YuvFZryLxmQzJCriMF309sAkRt8Ps78yMSyIZBB3xp6YK07BELZ8xIl4hW/ckjtW+9SinJ2tDCgp
l8d1O/tbF2GT6u4+DQOjszeKHSFyBGsrQvTnjB4QQJAdrtPR4NovW4s+yPQvgTtDqx4GmxEIqxgY
UKILAOh2xqeEbeV40F+Q1na6cvFSIVPWivpPJEZnJaxziSEBXBLGiA1PpqApDfln2KkKPb2q36kf
tbdIa8imHxV9XBxFNPt/aB94tKW40Te5hBfuKENAq5+tPgIGNWVQTFwLTQ1rbRgFEOq+FbP8wOao
hcH7q+KJ5/RDH+KDfTiCitRMtARp2lHLL6X65dy3+WkesS0HB9kJKsrX/jmGjK2FMawUo/jv1ErJ
UMRlHc9JgEEmGNdqNJpYPodsNkhzBTFPY7BfBg2tqEfSCcRuoMYHspspFxGlIagyWoGuda600Fsk
lXgJXL5uZKYG21SjN/zlS2FtgqGPp0b91jS/G9IU5+7fmUbdvRLz6lNR3iaf2EBYjbyczmpdXVgR
DYevP6LLHXpZA6MdTZMzzAHzMSvBb8c23XcB3OeG1Xh6DE8S9zSfUDjjhhPOEx5LSZN4qaJdX+tJ
Mu9UeSv1ElyE8piyYtBDSiOn6MkDizLAy9c5KPJG3qjeNXmoACGnLhwgNuvyjPmNdDlnqTTKwpgq
5FUVm+bM2u28qGFr5+wl+5BI7MG7pCevy3atLhtAmNGel636xllBnvrKITxjqSX5dyLTaPEFm+YB
ddhFOKiSgD70NW7z1KHPHCeLea4dCrH3eC+3RiggFkFb/F9wkSH9Q7HJ4XJiRzkT5folGcdR0XsF
LP/CXzfc6XxpDTNpOyLyFS937fVnd2EAYDep4htRCu2DZ8a4xDmQyHEQ9Y8stawayB2nLFqI9CWJ
F/5jE1S4vFZVNCKMRHrAtXnp138V/bNBMwvNRCUb3b9v98f5EWElFyY9+Cb5A684nkDvHbdmgcsA
ZJwJF373mmSCJs/Qt02hsQhPFq3vwMsQhpNafTadwXRz4VCJbrJnJv5rP+8tSc7EeXgYUHAzsQ3w
GQ0O/mDSW6nclf/gPyBbRx/O28PwfS7n1JDHTv18xQnkKj7KH49jgt1YkvS76yGEmGn9VZye5ffI
DYEtT7QXbHthFKGC3FGVJkMiu1bN9fPGDRH8rZyVSUXm7/8/2WtoFHFChmDQ2dX7EJKaQPJSyztR
udm2USpJSkIBJ4lkI48PL9ey4ECBGqNeunejY8a9mfzYZYC53OEPdt9FP3cb7fTdo2cJEgjDSaU4
7cqnZw81493HhrBDrr4kGP//t4Rkqi1MoTRKl12nN44CMtftrAB+A3EgkQ+lL2huDcPhSdQbmp4h
88A2ocf2NczfUsugI1LsIK/D7yABflRkwodCKfEqiDp3k/uydMKaKIGdYT5HhGYT4q4V3Z/yi5+u
h8ZBf5+rNn+GDF2cthVdCNrrwnao+51XTNERSBjxPrp01uKZ9Zjs5A5wPGMMjc/uDLGhkHBX8CYX
QtuylLt+FGhVXm7IQZnxzLAovQ+D0pu/qGMdNfgfxknuzVTFilUelWWOP6Ki7PFNK0JeL1Ygjx+R
k5YFycq9weqMtFiZu+9L3Lp3XJnxDrOfXCBxtHbfsrIDBPQglIBTEhTJgOqb3YlZNWWoT0zBTLkZ
RtNk/e/f8KyvEJFaCwYTwo60e0kfWZ+buBg4jc2rLUmm6fa32dtlirixpYerm5PvcTO19Ve5NiQb
h5dSNEWDIZaKNDK2Pc6gSU9JamDrQmH0Py4CmMYqd6QVlrWBt8IyZImPOPIi09Vu9gZhwgIc1yiL
13NfYBN8ZQloHw9+Dg0kQrSBOkIZC65B4NMIQD+1DKdRY5y2jBwNBEzjonYIdxVWPTMk7lO4ZmR+
YQKrRsON1lSwXOhcXn5zehi1YvGJFbE2pCkKOrR28ViR/WxEgujfQnKqwUHW01b0eR4STaegBmEs
DDNtqApVOFKjti8TIcyBCQnaGPmzKJcV3MkRYdPblHdkJuOq3pCROA5+38Yw4JaAmqivkbVIQWc7
aKPQFZiIaeqPXszRlm8QeqtuAV0zx5KWm/oC5ZqC9b/6+6LuYgd0Gi751+Zpk0ryMSivldTKYFBi
9J8O/HydCUvBAAHIwx/X4LC/rlvBufYkDv/rsImWKJMCHQjZ1hb/185dtlx1DkqjDYCUBpG/h25N
V62eFD54duMLs0JrqqQR/Ln186T4OSRb9OpoiBAVLkuW6gg31bljCjhChIdz7ESrxGs+fHWfHcQR
B/V5GakKy5eUMMhAE1zEhlg1i+OqxenY+aQNQo+0AG4hrTUdWHcLU8LHKJaTEktN11+M5TgrVR/u
zj/abNFUZW5Ebz0NnxicR9JnmGYidm5HbYfzfOI4rC0Gk0syk4SkfbCt/b/OEBwksUjwnCtpRrDa
MOe/omqoZM0Ej+DAPYaybHSE95agh+S/J86afi3/oF6ePeRbrZ7sYDwKH0jgbsMUPExYyoM04KJ+
x+CsVh6n0gMuWFtcN4RWefb6XbCtHx3esxsL/3JRGxw39YQU9V+GpBclW1hRdA3Ek/V1552JncU8
Bh3whKTygIbYyOYfp/9+dQ72U00SqeKUyj3BIHxGGEZkNMkw3dHwkSubwUmSTsK0pxVVweQw50s/
A6LNY+z95cOK21NTKoiXMZ9iFtA+BXI4v4n7/hZHJT2E2PTJyqx4oaWdIeN9mjCTg8hweYQqaQjx
3oNEMGAUfGX3vEMcpFjTY19SldpusEAcNH6LroJY6cqh43A5XIjv4IjJNanRwvMUeT6bl2YZ9UmJ
oIliUbfGgVkLDrJxFu4RQqWxJ1r7KZa22OHto/tMWQs9nq2/S+DGWwMWquY8XiFJsxO+IDJPSlLk
uYXsCRRedgz9gpB+JFJNkG/rzQLfhbX6E6Z1P/eB0Wl4pgHb9w7HPZI1hzQH2h6E2HsB/yuf8HcV
XGSHPK7wEuYan22CsjQS5G1A2Vr98KvM37uUDU0qK4UQ9H9/64FRnVweILVR9bCgMORq8q9XRdrB
1Ko/yrWSVsci7nP/hNP9uT7QaQb5T3eOorK0v1VFxPCija3aIK4UQqz/z5+lrPU3gScogMTLK11K
f6WmeW3Y+IfLdJ0llvYI3gYd5X/ijv9dqpBs0pqJeyFnhDxQPIWhkoi3Oxat3t80v1vc8bis72Xi
J0j7+CcjNbAPEEwDszN9FNpYmyIhSoLGhffm+0c7tjqnYmPIyPnPC3xuN/leUrrfvWMHGhKwot1q
3I23oxhEvxXYMnm9/nz1cY31eDkFTF0DVOeNYWAFH44oxgrHqFRPI0RjrOpa29Ac71uWLHD/ILFz
NrN60NAsMc+Z+MJrYorSKLY/VmHQrReQU3Ba6EqSWmUDolP54nHhunDKnjljpzc4DqbhlpnPsmhk
ME5mQHvfczrP8mu2YOSt6VbaTyQ502AlPmtjpwHg3OysWTnOplE3fp0WwvloIau3nPolVBYnNDVG
IKTd0QINcul5ZLyTA/lc4va2+iNz29igbq2xQBsgBKvokU357TfP+x8EspIQ4oA9jrs/vcuh1Vs4
fcOqJJu7k8KH42d8O9HDukhZcppSRKkEbuJrlYclks/DOYAt4syi0BxzdhtD8U9RuWc1WuE6nF9e
ctw6BzHkDnAwOyL6fY3GcExcLVpmdR6a8UdndbpZmBA679oImDSpUwMGspNxywI9pXHoNQiOV53p
mQeqkRjeWRGB2EV5GWM7BppRUNBytuFaBaHMckoJGe11/aoS18hqTv80WW1jQYoorP5mANN9ioAR
VTbDL7Xye2jDQFB3vD/bT4S3rKg/Udln2dXZdSQ5zXqJI8Udbs3TGTM0B9Oin5UOV2axKn2uavHk
cZDQaUVehr19TxIsbt/17si42FR7zLSEEKefQx8gCs/cVzsFLYZGnZid+QbIMg4Wzmev6u1LqWno
mZ50pgcnYUsA9oj3evp0dauo6GcZt+skGiZ/0Q6qX45bSV7wVAc6NYnVIzaz8BkjQDpUwyea72ET
+cQknCsAuALn4rviEQgxOdcXtmCmWn3GzKIRMgnyjKmadz9vXUx6BqfazH1w7J68PPQg99qleUYn
qioGwje8BRNLiC1gEC8ch1X0ywZPbDfl8uTCoaBHiyfhLtVHVdQbSJsPCTZSjuuYrOZiVzWDS6PK
a7RY2jHm0t1/2yi3japECzu6DcYbAFqOv/ntD2r3UYvtsOjwGmQuJJgtcFLyc3mP3PVqZ3CaNWVZ
lrnPNlyIXnzZk3hPY+NUSZCfz4fE0K4cnwqkZoMVdbh8UdFvO9b+trc5W9njjUIipzTR6Ksbh7ms
dQ48fLnEBUQTG/oiJXw3VdlacBU9Id8ni8jjIiXqe1yEO6Qp4WSqqXmH3qOdK46L2EHHSDkHK5wp
FJnjKaayo3Y1cHNPxttWgdxpsfbLZbLk/Zmh6tXHGnbei6qtplH6fZffzAENQNKovrKtI3LeUf+N
86IAujXy0NRl3DjcmAAZKXybahe66/zg1GL+FgsvqPBFVpPOSGuctLHbYP9nQiHVxSdX+PBI2QHm
u3YXlsSZNtjWkCBIfx+w4FcDou+2QVoG4fjIgrwOZj0Ixs9cE+xoNHPQStvegAykPCKuhT60ziB5
iB4XeHVWt6GbExX2u/ksN6M8ghmysQjIjrnKHOD4qHQmanICQDmokXTVQ2W7sO37+UZaK1GqcFUv
mNxkpFQ2QfeCxNtpwmgbBAdxQzJ0IKZNWhV18uYI+xVJ4774AxG/aWUz5DQ42uxHxE4rRQmhHpQj
IvRMGzm7O/VEk0K9UNuJTZfUcvJrVpcVvdefnWJXkqjTB4VoyW4zR+tfs1kISjVqoAxzFW/1Q99o
N1R5LqQLE/fEyaepJBgSSXhLK8QmPhBvw5tJnBIUvstVVta9n+HcSL+g0zZyDKhi7lTn3YcBzBE5
SdIlTnwmoaP6wfP3ConzE5ee1naTW66xeA+o7MruN35ICOvX49r+qPN8MdEnQxvbRJ2OEwQR0Cs4
9N/4f1/M/OXNhqKkrz2ZCpVVJup4h9cRNQYgFdXfQuCrSYhrv1m0QbpvbCRo/u4vyomikU0yf5Lu
ZI8qXoLoiLAJ7KiQcfKHuX3TJJrn1VrmLKMgOY42nFSMoB9/qn8p0m4WQMV7DEj4w2oHpMnKMbbb
LudnAOYHoTt6t4SMiO/EzYdXUAjAC28HfXAWYEw7mZFvtI/EikFqaGPppmY8ZwsW7qDGt6pMR+RT
eMNXXjb+fyYc6DAbuugOtHjYXTFg7LGuMV5J2YrgdjVVSuS40NgvAooL86WiWumy8GllNJ4XPIzE
jzjcBq1KsJ6ZtEHJI0SRCBO4dGtM3W/hhp6GoyERnQdm+1+DL1k2+2FeliKseIkw7jGagH9bcofI
VghE5VFAcLnB3ApHxfWzMdQqQrqoMDfoQv+v4icj4VTFYTfhlhVPZ5ziJLaRoR2mTxEOL5AkGRmm
rt1O25BwL1Rt1PhsjWZqMzAJSE1O3d37p7fOhL0bmGzfSQ+jOvXobi5t4Z+V92RRo/WjUdO+D350
urDRyPl6LyUabUcAbfsRQfajCjvhps0mVklK+Shyps9PQDBGN3SYkvO5ZZqUv2Dxa1XNPZp7/x7j
yLKZzRLwe9Rp5hzQ7fNuZWFBfxeKPkSaWMNe8vJD7cZamihVosKopTCbCIRWLhbF+ZPA849FBvuk
ytxn9xdD/gtZY2LJZ4GRUyjBnwdXlP6Axvx9Afi8sFvjxsgbER3GCmpyKL4wk6MfUfGAb3JaEKd9
GN94fPLGTjjEIbEKoA6X3y7P974zi1jJ/DfNbOGV62wR4CZVM4b8nAIP0moJuE5DemHQp0Dko+AP
nf5y8NY8bhs/QTR86oAb+IfK+dIRsHJ+cHJUqSBMtDU5Sr1lCfGS5xjdzFBQ9Ga+0ez659lFTRpz
4F2PqEyaBe6Q33QqAw7UMIbv3upOcYwc/np+FpPKKYCSo621ver8fLWBgRmdrO/9hkTEWcbEbDEq
5dYFTN6TvNVwqp+gOthRbCyL2Vlk+kMw/2hEwpSZOQz7xLq7WTSzHHl7kQaAq4ED4M2pEerQu0Ko
UAsoZFANTiQZLJEQZks54gA6pB1ibE7yK+Q7I4NMEot3UxUhqobczpmj3kiwA2WrrSqTAOBRku7W
wzN+Gcz6In36G7dtw5OrdcJHi2qw25ZX8IZLJSXdIrz57I1LRZQOgh7iG8K889FERiiMPfMkRKuB
i/ocDGFbZd7k3pU34xWJqszzk6IsbY0NwhiJnJQEYS9pgXyjjubxuFXDggjPkL0GRgANzYBQcSjI
g+xsiEQGSYUN1xt/f6lufxp/qVR2Udj66mL53RTi+zGBGNdoNtsVAg6E/uuZ3KUrWb6Ka3nbgwVp
FBARV+I+oesAAl2xPx713anMxIPqBHWvPorPPxdd9IQOM3oPofXjMm4NeO6xU266Z9u+W/vJWeuL
M0lglQzzdqEWKzMApnE+ViGlKVlhCT67KnFZVMs5rsJBvysSANa4f2dswRG0qMGvXYW990S+qdU9
s2rK1crkC/Dv9C+VhQwl1uRqedTBZ44qPP00z5c9FRf1712mGqRBto3CVVpo+3kHKC9LwqHqIeIi
lm+vLWfchH1aOxvRpKK1If3vTX2cC0FF0FOSgqmxDDqNptHCDEv7Xtbm0dIRLxmylTj+XPnK1yLz
Rnss6OR+/UZ2EK5EgRnGG5wIGUhZsUxRjaTN6FAt7CAhSg31/exgTalEds6EH5TQMNuFu/Y/2jWs
bdN8/+VOovQQh6HwFJJokEKLqNn+npYfPOwdBlZMA+oLEhPdjoRJVA9Muyi8yCo7UzYvkTa1k3YU
Egn3Uqan+McgDjYR2hS8kltY80Qjo6ZGhoJ+FaNDplxfDQFc70Fo4yuSn33w9ol8WjXovlDoGBCk
LGmYowwFHJHQ2Iuxgg7hWEj4CJt9rKc4cpuZ1lzCoWG3mNn+/qtf49IqWIeV84EZaO52bi/TJWcx
CXCivdgrYQ89EXm8CmTdLrHYpqiQTY8kCU0jZ3kWpkLORW3VBRkKHlcBUEzLa+svbCNFGVHNMiTi
q/ZmhfI96SHXZHIlJaAQMDV4g7rXE5WKr+fiJs3NyeTap0GaHfpptPu1EqufDHYgpBZBDZmHL41E
NNR7rjNYAbUFYScGx/UDJXzboUMfzKOwSQ8b001H6FpH3KSHuJw2D9K7AABZBDHx68qvj+obIAmT
eATs5BkahYXVNaQxfSL7CbmXuNuKnmHXhJqQNvegVQo3FHQUFPKDRl3i8P/8OrOwvLorJ9xF5tSI
utcT8JIt8itleaC5acaQJvTKTWYEFMSynkyMKgtKYp5WcuIqPtxqtYlJCIH15fqp6LDCw4QlITYL
N7xFBWhOBlAzRdiVW4LmC0In530ETHTd+pAISIUCz9MS51nvE6xucktQ7jIQWgQTgo/GCGvue+qJ
bYmVK6QOYhM0j+TFb6NRHNX7HFKivWiZ7S636FlPW75QHbmvT40QMxvR+Qh7yV3m7vCFy0BPZdMq
QTrAhc7ibJ401u72eWgkTUw5BvFeWdtoIbDljH/VPdFqlGUeiwz4GEh/pVFQj7NdFwJQqu853ddj
iLIpV7mGLMnf7xyj/iOp1M0IIbBDQRa7H661W5C3A0ENrn7MazgU8IcWpJsvY1HwhyhyRH030IvG
fZq41KCuIGXS1ckxvC3qfpSWAp7mjIDTX7QYonnHd9C4vPYxEQKQPOqsaVAyNXwpZ3kX1ccH8cnJ
ysGT8ptinPcK2qKrYwxtqY1/EQcIi7O6pvpqKWm8TLxkiR19wukXN7cpQz+MxA/ZgCOu+oEk7KO5
sxM5QqdTZulxmWYm1blNNS2FL/GFqkAeVZkVrIqCdiKqWrCYcR3QFjHSc5PEbUzaePpCsSWnwDtp
hu+C8MYxjsu2IAg/i+Zk6FMu0YrVefIY4A1A+Mr2FWSqU9SG5R9clRDbjhDYNYC0YRXUkNOFVBSb
ypB4hMoNHCBh4y1M036iTsH56zeH8VfnU+8nst5n1nTcM4OrLi8M4OHTCMtIAs4XhilEari1Vzga
Qm+Fo7B88WihRjZ2parSrk6Ssa9FjUizSn7hokuHHw/cSrCSDwvvqExXBfKFxQxQt6E/lDyL5VI9
pQ4g/g1+4EjAdLUrd8j9xaGG0peipRkUi1nhOhHBsYfyzZzHmWcrkeYvDf5h/3K3y6dT5t3P+AiX
147IarnxsPVc8Y+5//QZ94kfMlSV1JA3qhK73p182Thqg8PVIRNVEsvMXM5stfCLGSWorNEnc+uC
a5jItmnv60vz3TfP3yAkSc/z/s+hWoZVjarMh9lNVuaQJQmKU8T5A94hZopegTzaAmsdHn87Rdku
zzPXzrejmKJTSPJ/QHYjw88nPUBAJMsN+Gvy7cVXe5e1l6ZNd3UbGuB6Ojnza2WeImJMsJcKo7lh
7HFQ1TTCeEENVLvEE3FF89VgCXbPn79wFXiBqKkZVP9IaRie8zVAjmr2jqBXh7c0HO/QA+vsPST4
os0PkxATiR0OCstY74sh0zeUK8aMKXhistnVJWw9uAskyyM/pMauCmLKCLr+QlKwT1L9PLtgUSLQ
ofkA0S+ymEO7yVqCOOX3SlFFburCKxVjPae1xEKdi9WMO0zNfE4FTfu5woS+oHZgJ0STt8TVxaum
nTsdlRrQW3rl901NScA0UtJKuhD4T0jyTe9QjgaW1/4QcDVsA7NkISQBsBX4fiEsyrGTZOQFEw8K
dNR0SLrKUKm5/id45Kpc0d0vyzznxk+U9UnMvT4DJRjd/hrXrO55iIqxBWpSguZdoezdmzuLtWgG
mcxih+2+Z6MhHWjSNl0znufRoMfNGvVA+b0d0rm4AmSa26wrlnvH16/eHu+C77FKzsi/Z40dg5Up
p3TDEGrhzrn374uKkB3CRGLp6IkMyQBUUp4YXrpn+7zOU5suBBroV6MmH9kYvoJzBwuJpIwAo/2d
0UdUzjpyNzhxr2qNebRhhUrMTjmiTwXPBtblOl52iCIg8dngRmOskNkDYuyis8bXapEG1OqTdTzz
PE5BryQCIXo+MTSGIW6blwUwYc8blFXE3p/e4XQ0AL8BjHfs6YZ+WGQYrtSMIiXwS6kLyKhzt7M+
3BH/0bTY2mn2Vs0f+AjAfdpLxMyPYQUONXYg0HPLAvt1rbOMz3YQxmnxEkGzyUg7bG4DIvEcZvLr
ZhWrYsXTVJHtaqaFcH5xm8wu8py6HHFKXNixCknUWhLLvEsEkVgq8OpXRkCbGvgGWlRCdvo4ItIg
+cRpSG24icD3JOzNcrhZkVx2d4kr+Y+JR/3vxIlPTtCYB3g1ZXDz5S5yez6y9qFiS74Prz1ghbel
LOlv5TQ3ckSZvp5PCRskTnIGMGqyrclO34+tUe5kuzB0Ksn61oWb3SmIz2g9Q3sJtJ633fy/gY1l
5LyiRieFhflhR+8upFImV/ZNDWdM+aBdbCTxEnOC8F9yrSTgHXVJxS+IE5MJ9/M9OZsH6aVhTIjA
gdOAtgO08nOAPVuW1S41yoWIQwG4vmpn9rFKosjpJb2jCGSU5qh1tOwQN2kBbsITlr87dDwcLqmN
aWy9ZCdDqj1J9IuLohYIuyE03hlxjsg69PWUF1x35CBLStDJU98Y+ofHA/SRHdZNx5P80Oju46oj
ye+X99AD2n+6nTEhw3pffvM+z5fOY1nPoBaIWXYczVyMbaYyAOZR0psn+4M0JGFPJp36XNinyYAB
44dzV9VaLmrxySfZVas1gKcABOQ5ECY89w1wZjh2egAxCoFIWTSSnFzZSE+chY7p+i0NlT7Oe5G5
5SyJ0fkRnT8h0hGHhiwoBGH3ZGzC8xDCoIduhl0Wmddrug1GU5VBMbsHkeA/6eaP9Ivshklf47Hl
f/kEwkARh+BDIzrY7kbGYC4KTMxbZNlLCKOdHjY5EeKXx9oPEnuleSIrivZTKteAIbLMUohCZoWg
d8XHD6jjImWPnHZi1ZAd2KGHZ+ki1D8jOsgI6a0Bo9RJ6h0Emlzpu1hfn3OEMBh8KOm7ezTX/wtc
Vgvtfmk3uFCf0e49mX4CXQ10lLwSjVO1f50zl0RheCEga1u/2UwmIg4Nfgwmmoflqoz4+SAOP2z1
s1D9IDUqFriPsSIVAY1tkBSeMRpcreijHnoYOFNTJAryjeS9cd5m6VCHPutPWWzy7k90WGt1EoOX
z0Zk8MZZFbrf9ctyRBLurZ6Gjp+Xc+E+FdSFVgqjyo/XifQgsHCz0LqNOM1A64kk5M8pjeqOn7xb
GDHDkaeD/dkE4K5QaOeNu93hhK8i4FuKhi3J3fwb27O7ZAoHtgHZNYUgjzxSGnR5nI/KlxNuzcGr
HQiG+ZfRE0PE3AiykfT3UtogHOSAg+4r95ovIycI67d3p9E6wbYlgrx8yW5x0gmsChzEq2DJWe74
xyIEIIGr3qUQqtQdMP0VuBO5v93OrTxBRpVnR/kJZL8V6gHZXt4v1/quUJcLjyd4gAXCF+RqcsNh
Z/ZTuYSvb4VJ2MS5xXuP8yD3vLof+pOs3K/srj9eQWp1qboRsRcXtZDTByOwRo36H0APTnQ4zvWM
pw8NWECvV6opS0kv2sQLwiXrbqUpz7ufJsDQ0stTFwUgjqw5PgQ3MSel2lVciNQL5asd0mgMOUAP
eSUwrjFhdbshSBv7YrTRInFuHhjdgrecFvCS+ikUum2PSXkLU3L88kYhBHP1P/jWnBhiE9L+EFMZ
JdmNA2upTkIMKHJMAw6XmgBy0YXhnExWM1ngzHYXDad0Na2OLiPMVLT9ggn6dTYwRZ/FtBvHJJfN
tCYc1vpzh/i63+Ao8r8aLITQRvUH+Jpi2cLRh9S1d7lHCXxuLe4DtsJ1XnkrMWHOFt0qSep9CH2w
bvLn1L+DaBLYdMy0npwMX5msfHKYAgYOaUxoAIXXc0tIZr0Lw/B0vgUMIvAcBT0J/zGe1cxhdCs3
0AuE/fG7xNJY/oC8radWmRY09D6TRuITFnVWTore2BVB07u75f95HRXwjnsmov8+F6xiCOhU98J4
T8OBAObi5YchXhnNl4YeWb8pdaMWoxsA90HnbRqzYZCnmVMSdPNIU0mEZ2dKgelcVjsb+eORv3Dr
18YSPJ5T2T+3UbmDjk8Vi41VUI0fIrSyA8RH1A7dpOzQ80+gZBeD8UEbwekuFOBtL/z101nGZxmb
5bl+cjqygEG8D9+oSH5EfFcNzjjLj4W9vtTQcW5GuyTzNIIzwhP9z30Z7My1EO9FO5dFjrO1FtXP
5vJzXuej4JAIUoNndjJWTxFTj4xu07Eczm88r7jlI+Zjue+r6XhgoIxW4iUnSX1l6alAC6cCb4iU
okaGUbzkf0Yd8JZcqo2j/Fndq3xZOg7KhFVjpdE9/pcpxGkOmgyavQhx0SpCUK3A/9erPs4VyihG
uQtm2n9IF/sPS2rqKzhBNU9hiuJzp3wGWtPhDA9UW2a/Hd6a+TauA9TJezz+e0W1sgO0CFoCf/Gc
Nf+4q0koZ9K8rsn51L1jLKlyzlrH6pzpv2c2Hnw6xUkED0KA2cNsouZb2LCdFlzmpP+xHRS3DSiH
EvkXDsqkdD+FMJf3leuuFBSPEYoLiViqCvnP5EXCnQm/flm8cohV2YgOx3Ys98ai8bMeBNHDSzvD
rPurcxWGSrQMSYjK/66w9fUWnOfyLMyXON1BHQj1gmED0nZwR/So7uOya+0u/pRrSRFSH2VHlPDL
CN/5OX0IQZViCp2rmJtmmCMtaB6BYEi4XBKKyeAzeJq2nMh84twL39OTQ7bum4Xl+9S1NGDm3OTK
nahz9A8o7vaqFweBwylCUDc53oFMgkOqnFVYN39ohfkTdVC7mVF8dmC+Sn4dtJbgfKk8vhyvmskd
sfa68fzh9CNr7Vy5sWgNhoC7cy6UpBU1udTNbdSbvja5RS31BwAJpnIqL4wSqliS1Sdkyk6vQte7
0YMW1ERRMj4XoOoc04yswnUa3bXa8kJGdBCweVILNkxpL1xEGyVC6fdTcJ6DOqLKPXTN99CS2cOM
NsauvTGeHjno5Kd4jJyKjmlVgpZVDh6odLdzkKOSeO0b8ZI4fGurA34e6ZcCejRDYh56qCxQ3hFg
CoLGDR6IPU9F981lOLxNj+4zyio2uf1Y2ShKUEktiBgnz5nz8+8h/t20lPE7pD/3A7BxkAjKLjr0
5z5FWjV5s5F7xRr+Nx0Chl2apE4UkwumFfscT5EVmy1Ll8H5dsj5HlmmvQqhYGzTmofxUcyCGc5c
tENyI33q8bYWD1eSAluaLsPWIl/A66Yvb7CITV0OUDjH3TFVUfqLe4baVvxHgfSdfIcfrecK7LXW
to6cpCevucY6jRgZOMeh5s5eRiqMf8jR0nuzJO0SAIGUWfVfpnl98hawNrbLyNei4qx59Ft/DWTw
TlNMDMkFCL88AEVbbROt0kGwnPoUdnLUcEGp/gLqd/z2R3ZzkwGR6Z6fxbQ6+zzT98+qRsZ+bfsC
yfElPL7xVHmfrkNq5qSQPHFnRoXs/2TN6cYVtsJKAaG5ihBXDrWgWrvWS2+vYi3t8ygyf1K+sU9F
Nb4LCMWn236RD4B64kL1PRMsw8ijcCNW5W5+KqlZ/ILEWSO3FtR8zF8FruJmZk3lenIilG0tqRTV
KEAyWgQOcxtg6AmiVlfvq2R6f9geXmPHsdBg5lr4r4T3b3j1lwbzrMSDWQdTPmTYHDr+TUG9A6gY
HA5nGU8OJueFPoTLjHFHBL5Tlf+C9nld2oja6zDO0+iK7HC7wn9OyCAbHWcbC54+L+C7zH0ScYId
9pVAmSkyK9b111omgV+gh/BvkWahvy8bF0sZBPN9wsW/Ikldrg0h5dCuM66Fy0UVKzoROdS30oRd
Rh1xILl4bHnEe3KPZjenpYIZGft09MvtU8y9G0UvBD4GjRqIR173ljonBzystu1kF384KpuLXXrP
N6gOed7REQGenYTWh9m35nF+s+tCcbrWB8VMrxBNKifKRXJNTGRQ3n81JldG93zt0mLy04dOdsFS
5Mw6ja4OgbIYC540NQQZw2TnSYgehym4lobYtLtM1yHSVX5On7f4uWF7TQUD3K39FrVq066GjMcE
VaJJeFbQUFZIbjo/z0xC+Hvxy6CkbaOY0uLU/DeGDuoYAK9JgzaUJNEJ6TwKIDhan2qo6HE15LaQ
+aTytOsnb8DHAZgdRx7HlVsCI3PucQcN4Z9QXMIQkOjQIYn29TN6+EolnouD+ynQ0I0CUoTRNMDu
Nsv9FLvxXZGr6YbWvz/XLhq6OxaACkPGFbzzEtmnOq9qc8FK+4eAuk4IWXbMYxReLOX3WoPQHq+t
Spn2RYuDyiYreqP6ALEs/yuzgOd+zT1dBPfs/YCuvWjo5wScrVT5QnBmEV/hkue2eUVqvqYzi9Uq
aU1nJoEOmiiGvFDo7oZMHSbwLaKL9EG0TuiUcURQGxnqyaNOhDbd2dEvmQd6tSNLW94S4vATZ3Dg
OMYpXWJt6qHY90VwfkIGs7EeFR7cdylAAg6xNR+cMHik/W4Gh3jqn1N5uinf/6eCcBnp4CzoVH0Z
IksZL/0+iytoY98RiCBDpxRRlX5cyrgKezTvfT8v+l6anxvhabbDGWHZ9gVnAoqAT90UfNuPMLXR
A04LvHkJJ9lW/eClhxAwmOqENCw3cTWUHTVJyOhXmCt82jxWTnVZ9jshjL/TRqgGYLEeHlfOsjqe
pc+feS910uBISbJKfw4c4kL+AfiJ8ZBeZb6I7TESpV9rf/BRhu1JSLboZVyEgBmoDkXKT0Kthaav
euCnPbW5Crx45ogL7n16EjHTUORH1JReVwAZTjob2b2cCrgc6bCMhz07+64y/wAPRFTniGhXnmgC
hM8WmPzBSkmY3jTeNTyY1M2RM+0oSsAp0BZLEqKA43P+Xk4Wjp/wJe1WGhCeg5gpwwFME11sokhM
58t/Wr8zmEQ3RrUnrZ9mKm4q5XTXtuLGgSLtWepgnzOckH9ksbS8y2Z8zA03BUZC9JxolvSxULtf
kaoUowwQ0pnh9X77vzOFKJZi0vuI5e/sJ/gflnzW4E3gk077XnEdf2yLf2Xgn6flKMt4Chia1/8v
kT/eratuKq3RKgY7FfJPbVyAS9Ks5OBRaIS3ANxf7/fHOn4WcMsU7QdvbokNlWCVEbyxT3vJqUZp
/ewi2XFaPLgI0pED32i7pHkYKHRYNykxjZtMwtEdlDoD7y1e44j/OyemSHp6lMyCm5Nsx3gbArv5
nnjgbY9zunEPR47shKUt9KGzjLYrHCuX274Bj5xGN1vH1QsA07bYwLXAD8Hx3pAlfoFwf8bAzPJp
tPUacE59IV7oWYAT0i/znUqzV+On9UENz3Hwl61XCyjHPWXj4y9ev5XgtrlCG7fT0zmnTvrcTwwI
1rpx6fqVibQVxnpv6XieiOV1CCdJrSnzyEvJmgpbMh97qN0sYMfi8WyCdP+1dZ4YMDn/2S9O1UTv
N63GA6KcKF1w9o6l2apkFUZpwlM6uvqIh6NC9Qvkvo5XYKpXcOlfVFGmXBqlJ8POa4CwBW8zJbBl
benFvjBt60Od2+vdAw96uXthjq0aweYLNRGNMAoitZMvMA7jpPljmNJkEO6k5FiSLBskOX3bMM7f
0pDqiWC6lVlafYi24QD2/0WOS2m1dQizEeHY/m96zarFNlF4+Eoh5yl/c4GluCrmy1pCJDC7vTux
cE9356fzbnA3JIOe0uzNFGG7J/YzxwRm2LVQmRJ5rH1w856bx2e7ek0phdP+Kpo4FE82qSjBgwLh
Qj7H8awcuTWJOcJEG2K5kJpzX2wsr8tJF5xjZxPP+u+RL6xDQtu6xHbnJtLhJWDpQJ2cohMdgPC2
WyHVFIeL2GgXlqrO3yK4mLaG1dc5BG+v7sA2lAK4Oag1WIDoShiE3G7Zw4qHpBeq6B7j6tpMy5UO
/cVyGiHkaY1arGNp3vMwy8BV0kEe/83COl188nA4GJ0bmNZfqXuy4h+gk6hu8L/b2ZX7ib8cWas2
/X7L0ohB/XCm29JHn5gvJwTBSOp3UfbXIVSMdWNDjgdv15FOEW9A4SKtfpS+uSJm4KdhgnDXXw5K
62mDEkEXuP+S5C4D4gyh74x7+rEr7DhpDO9YAYps/qSdWIx4YIPAp/8OuptUd+3WzPmlds9EgMzl
thQFNyl5x5Tcpb/YuKPr9ptZ0onR1zPuQ/urjaVrWMErxoWfwvuLue0JTjFqiyw22a7PRTrCnDLk
A2NRnCwykn7PdLqV76Yci+1siXXNBRUFyMJY4euSq5yQkzVHbEYZ1Dj0hBcMJSQ3pQbBP6eW2wsY
+UEJHhK6E9JwuyEbHA0YEJBYCUHeYAbNcAM0dk91mygRsGKYucFfnM6UaBmDfzxJWrWmS+gRiFNa
vuUmqVGvcRneFpSjbBxDSCM5mvAUW/+rQv0hR3Ao1N+iCJ5yKX6LuQxb+oHjAKL99RwZZm3XwLab
rmwOrOzYWEI5lTQajKcTnyZNaCT4lCD3wyWjOpAbu9F885Y58Vi+61y0l8NaDWJwG/SK2Qgd2KO3
ynuU8Vq6n53bMYz9S5LgnTznFDAHfBQETIzhixeEu4gXeM4b/ldJDt+7eKti5tvvVR7HX0Z9KOXP
fYCBC0CFfB4MCi/2r1VWRvaDgrdWoyxix9IiTgy8akCRNTBDbqI6nwLgh8Xs2ZxRWl2j4EMT6CGe
DV1wa2xjHm9uGrCYuR1vFQqSOTGXdT//DxsEDk6x1mUSsB1tUFcnnf1akklFXWKjULBzW0GYtHbB
GClWR+iT0Y6oVUeL90cd7EbQw41b+I809wvT3i0/J0W0i+iRn1CZvM4VoUYva3IQXR/Q5FoN1Tah
ateh/RcBI0YSFx01noR2g+8xqoQA53hJB5YPi/552AN/Nb572fdQE1j50rhr0XU89aE0dUdOIkX6
e6Ex8pgpjJIiDZJxZmoAb2s6m8gJpOktdjQxcSFDiSqlEtrJLuLyzPcMUrprADpiaCRqBYtzkxmB
a8wJNYC8iVq8hxGLQ1n8HIiw80sHzUuRbarbuRrHhhc8YUArlLP9UrbuqZizPyDwHsea/FgB9o7m
ifwNLoTSTP4OW3B0YzS4kkaq8VAwnsXVrZCaSlmnhW1BuIAPtDJOabWXpwPh9a+VQhMnNfjv/Auw
AYV29+iDZOqbau3UcbkpVNr48rCtUGZf5NFT1QVz+lY3rXIkbKgDNVmixUGwF8eKEthLJAloIeUm
d+QVJ+Q1u8gBU1sDCb/GSvQntJVn7uPq0rmUQbFSoNacdBPMFpUT7OkgfnYdMQgWTCgIbUJ3Nupz
2/dIdrX3zARTenMH2zQ00k60Wb8VJRtmb3EH7jnazS38qoSnrtYDCwK47SlFVXyhSKOZjkf4MfCX
K4CdvtFxIDE4T1UtFoT6sB4BWilAFxpv9HNHV7pxH9NDUTvYp0iRguROt8845apChFH/zegwDftP
ZDAPS79FmrNU57LiIwljO/wrHVy0v/7TX2yb+/YP/ie1mRIYljfnWWk0GNoAU7YCE89AWdzYM+fv
FCNaYEP54NY/5Mjn7iO04Ux6X3dI9R0qn79Vwiy/SXYRZhneoVYgrt7kSIS7kZBngyoQbeW+KNDM
BHflWyfry3pO40DRdp/xNQPj+ofjXAgIgHF/OJL8UDoXFTnQd4La6Dqbdzdsdrf0p6ij481sVrAU
kKiXlSng4a3xYMmLyYW6wcGgxBJ57pgE50C5NmO0OFfS5zDMsuBz+CZBTuuocdobV5WG7ud7DO1D
Gc4o3Zbq5D38zpsSn9EwhB8rEdVs18yQpTw2MLmJGtqZN55K/2xxDWeNOP93+/z1GJrGkMw2C8AH
FRkFfpq8rWuZd+46KTkI4BJycTnyBZEc3ss435+MmmuKs5gMDDZA+V9jozticnOKgVtR7JziGKGd
vV/ns+6rrioHesi+vLXdiY48Y3kPdLHqgFWZc2aVfk40SVECRFYj0V8BMnDWSdQo+hiZADpCcUx6
FWMren7sr1Sov3nAKocdZxWH81UOLrASr3kJTWjPHOV9R8SZocbmXXLrNXp2s9Fld4eygaDtm7wd
mGsoQ4L6woWZTTQ/fEpFRlzMtFo5UTZeDeXUGQfTwjFRVmUeMjlktjb6lR2gyfUij5Jw4gZ9D2FH
y6DWIHJ+2nBqxSVeIV/nSlh2Nt1MNOshqY9IGVy+TU9zYqnu776FDNbxmUgtPlgyqiUyyGudi2ox
JubVfYOOnGcR6jz78RQxpGiBUtV7nkrD0XhhII5C0vDuyrUygrf8s61T9aSIcGBfPmf+N54nu2Ms
Z/R/PuKAp58LmileaIygy2gsrfhuae/tfbKMPX5ZyYTu7O4LgnNAym5WYdUidgjQ7ZNso/1aeUkU
Y+JKl06xXs76bBcpFyMjkIHx3X3fybF6KnTFGafWaeZ+eH396Q+bZlNSJ8b/oycCM68AUS4XJ4iO
AEf6iLqoGex8OSUeKK41drCH3Pcm3mxAnBHb3IZnTVuB/BO14Wu2BTuSaykjT4arOuvUdVnz+Zh5
66QBejBbAB7QoJa7ofxyzLkHVjn3YgokszPw3YepdWduTs2GEd5k9tw7mckDZGOJ2dNI78VpgW8y
zWodXMNNMAUY0v3HWr8nIfNuSoyqHaN/iuaCt3Vz9uO0RFoATTWKn+IGpJGLMp2ffoFFIikBJ6cr
o7860OuroCmY61jKdyo36cJnskswOB6caI9JoGFJPadUpVtEkGZ3tBf+BZZ0CTJ0LdWc8lGmxYOK
UssfyHF+1vfd4ILDhU/kI0SfIPxGlDqCK+xvTqtppevxJV5MZpi4Kg7FY02IJNZtEg2onbTcxv4T
Pk1/WdXYxjY7FafaOCf2XAh4o10t9Aw3BnmDUCdTQFa7GU0aiOKytUlRVNuTvI6qyxDG8NuIlNNZ
mNcxyCTOvXp3c8DVPz/Hq+hUj47wqIisd0NMbwiyZK7eikEHjdBGvDvZMRNioKtxalj5LrN/cUYW
9nJHKOH5v8HZlMtZHh+ic21cdtNcql2Aqdodq034DtYi72tVpt0vpty0Zarnb417ETmbH7b0DsKl
ofsdgS3Gj15bTaw+g9SFJ710FWyqYl4fF6Lp3Mvt07DV+MAB/VG0h1SjXJmjkdUaj/Wfh0gmI9zI
EwQ2bB/VwnsV15Qn/sGllu2P0cI6vCvG0VmyiRUaTlPexAfStLgbNnFQsrVqycMnXyx1/jJg8R19
cR4eV4e/LcT2KsNL6a/ZlcT7NFAMoFQSmLABuvpsD7YLi9r+euD0oExuF2amsf9JROtD4W6MsTkd
NEFUrOMxkBJR4dOOQwQmABspHLnVfXjxhGf0EKDXNSObDUAET+cAby9JAxzar9ARtqg7bn2/Vbu5
EMMYOPSpq6LGnNTesLML5W/pEhC9EUq3685+S9QMMwmKAErG2Tdu6xuiDltJvnV87i5dZWlb4T9t
HWDvLoKgRRQ00PbRTNOQJU44n1YcY3CtU9jXI8UIMojgV9TMypUXJ+QhEv/gjxIm5C6rTAvY0cPa
PSLKuw34tbd74jT/mrV3CZinEUQVLoad2ETrvsS6VgT+8x13sgkUt26cuacn364mZQ8HmCoN3qgi
7SFZwA+z70tgRYG8ObNqQa/Y3RjKUnr05emDxW7qDBFwKbgsYGXwqFvFlvzipWTYUB9KgL3gDnov
ndTq7Tv527pKOCZjVoh43pkiKM0XuDXuhOFvfrT7MJe9xLY49lEVdgaKbyobUE2eaAJqWd3mbrxT
QOwlQKdh3TurgQ6rLLEMunysYv0Qc6/ZF6Mjwcui2F/PJGCunNNzr+Y3KdRnnsLD+fC6Wde7/Yaw
XW0ZdSrXF4/+ydiaBxGctNiOdRD1CuTr9GEVtZqldeDnZ4O9d3r7PkL/QPhILVqd2tJKNzK9Eke6
LZyaYSwKR4cF3IIen2nUSxGlsAtGc6CNml//ZTCZw/Cq3Rqtu0w+o++9QaCatYAMXUsBJjduW4za
PNbgzqq9M1kvcvYm8R0BpNnR/vBncpLkaYQ5jLGEMKqsnKG21wR/roUhxK0vEKKJ1xCzQI8Z5hcg
SIVbNXwTN4+OW1Kd6sviugWoDaIwihdknPb3AoiNO+AxFzZF+tVCdORfKVTTXglxiLbndOnm3OlL
/wHhD9pQdcE8hgcFuy7F+NbUvYpWl/58fVhY0CbEzp/xAn5+MSWRlJagMQlkikru9GpdQgDW4tRF
MkWBB6QSmz4y9q6IgA6ddBnNq7vDXPJuo1MfE4QsJuuFJBWxt1DK7F0wpkKBh57dnzOXy/jLrAxj
hJkWhECp1pvv+LhX3gv4oyZsNv6FDfMeCzLkRarbpqA3r7966/ZPopYE85a42V9RA2oUUGzZ0FEn
vaHwcvV4tUGC7nqYux2aPJKwPEVn1vKQrCASGB+47c89DoWlWiY5FdB0YpkjWbMdVaKYKUs6MiGk
gUZBkWrtugJmUCuPsla9rNuwnw5Mfe0rQKSyd2SI2cpzo9PRjc+i0NGzL7CrFwRtGau75mKcOXRH
NlDQGfKcvXMBpSJ3xkwFZimpu0p89udDunA2yPIhXUBxs9xodwCaETDqwOdH2bJlUDNDdT9Z8hat
chCeJJapAe5BxvwSNF/I5dXfF3tLjWvwpxcLwW+xgeGKSxnozdU5Az0pkqcDg+Xw9mKXI30yr9xo
7+wffnlbkQxcy8ZFB+knTzFPkc/llrvWFHeEh3xVN/nPhKJVphvZeVPx0SlpA8LZTPkejK1vfN+o
9T3XIfHgTXVfwcYLGXILYpkt68blSmmztYtLK+MYFf/EuF91rfV0V0ND8yxC9ouSuwCKDLPGpYfQ
Q5H8TNdHIU9TVRTZRrbcpRWieokzw7dQDi8hAyR57Q4PTlVsjib8GAxHLcOZcEvG1+4OWoEzvZg0
fPw0ZfFr3/4sm+i/5Js/aextBl0/TUGILUCMtDaXNjijkX6aIozqLec3LLwXBzRlVjbGouOLUQXS
PUkgmyJDC5wbnYIPzcFfPaUb2twCwCW4cU4XYEfrqv2HLuZox1VWvDnO42Blp597WLEJPs3zpvb+
qrlSD5CxvGDSomCqDrz04VBZOLfrHh6wZSMPejwYapDQdGqpzLMuzLPGjSoPors7g6mIyDJMcAwG
wnbTwz0mYtkUH49JfvA4bhgJMi3PQXt+s7Uee5vvnBT1D2avYfwCpoR3FD1k1w6s/KXxQJC+Dz2N
Dpgn25I2zWuxWTNFeeQLpjPTJCVhpocwt/N9MPRetw/VebSsaB9KSxo2GFo6TU0FACJ/umZ4gAbI
dXaqyWJCS+hK8qCyWMP8lCL7E4DUiyoh66YP90A23GY3jS/NJ5X2NAvNzSgCj0FYVYNbOD7br7r6
yZN7Z35QcwyKfyzDsluhqo4nsPXZoZgUGFEHUZfyscUJeHFNlYiZQjE/qkmeXZSOHs12HJmaH+fz
ErRNqWJkeKe81naz0Ie+GhaToRljHJIoSkAbec9P9hKlgPaKGhXg7o1AROZe9sivqY9JRvHG50GN
qQ/S5Nezq6z9LvOn9bF6D8zokLTsW5eJj7XEC2lec0vtU7g2U+0bQosXJlDPFiBKHqJRbDPJDj6k
CbFCEuHL6URJ5B89/2J/1r/+dcLyW5osn0k5PdNBVV4TqtmWcFATdozwReGKTVTiNiStGYQPFh2S
jS/Iq2I3+apdT9T9VnZHNblYBAc4jQCRKTysZjPz6uF/hrsrWAdX5H5RVJu6lO6o4mAsi6D2cUJz
Lzt85FdfKM8Yo87nL1UPZ2y8iAP0yjsqctqqH0xTTQvx0J38b2slzNbmbRPQj2VV4EmjX8tACGkW
nThlv/+wfQ/FKeRGJpISiSR58lCzOXfJDizItKdMdO5Wn99R9hxdfjZF4G5PypYKmlDQAqo0z0Vb
2C068Cd3Vxj3iQy39yf3c/im4P+5BhWFa25NATvdzvkwCy7VZdBOfqI3assHy4LmYxh5svrWjpmC
ieoal/61dZZmMG9WnWU2/TJg9k8t1LjoY3wkOW95YYKoP0jXWxEo7U5PhDSl21xlsG4JAsp0tiE2
aJs/UW1czLaO/Kjx3ZiEI30WqkIdEKy1FH3RZo9yQ4FPC3wuMCb/ufN3Y3JLyC3xD3RPdYYrzAXl
ziP0GR8dgsUB3gwd0jzBMkhR2M7Jx6/aS1UAkzNz0t6O4TwtetMo1PJZ3mMAzdQNU3TlKNnnsvc2
ST/8Cu74tqKSEOZW6LOsa0cAaCBk9PM9Aj9MJGy9YuPPvozbVLkDzg13swELuuOOBCartV3yQRhi
Y19ryNGsPl+vQedBLIUwyE3aFBfe2ihlLDA92HabjCbVXkH9b5WBfU7UuNLsnnp+4mux4d/bx0u/
4Qi7tTUkAaYGsS2EZckx5odJyjr9OcTE+PbkgAPZwkyh+k4XJlT/6sH7JzwyCztBWvT5mm/rpwTT
h7Dtr+1l9iwVOpGBYEXN2czjJm4WSaxcxWLY4aqYgZkxfhmozaTvhPM+jjtjfH2isAn3KDXAMKAO
eli4hFHJKB5nHuib6z3sbyUsfB4MNQiGJxHEnkKf3fNukz9VRRgH9R2T/fFdjH4LBuudjNa6sfD7
vXMYxdot9Bn10oNKNYJQvyZsrm8mwjlmnxZ6hnV1pgZDDhj4MJxVNLq5SCPSlJVgtru/RV7e0DM6
RKLR8NGYjS0V4DlotPnrEJUzVF1gYEhFuPVs97zKVnb81EYIMtUftDYYpTkPwDtWlFz6w8JDOWO5
g65QH1i8l2UwaYrVixgNYp8Gn6d+cQ+5eUxXl4qrm5G5p26lUUXt/Rzdi513v6XkZuV0I12Qxagt
ihID6Sg9q8PR9lFePxkJMPpHbNr5M9+/ksLPtrqYG5wS9KkiA4Cji1D8L++B3H+Lmpdhw+tbd2s9
xBONUpNE9hCh42pBriZJCKItlB1B7ePvfZPoO7e/BxFLQaKBlq/NIFkZZhHWUQc+tGB1qjWRm34z
YVBHLCq1BNrqZuHZfP1XJwk3AUVAf5mTrZL05swJxvYG9ONxrnwVTx2M/SNLgvYn7FscVq48uFot
4FWpJWuN5lZ8oN+VFnGwwuz+Dtrwm8L2YESqPKP9Cmn9YLGH8JdQICqslPqlg+4Ae/269icIxrb3
/rNS5/cbbYTQaVYH0srWGuVWfseVAFZrnsqyp5JPDFoq5eBo21p1PQA1LJmbfNKD1ynpjkwfC3LO
ZA90RBQcs+mgxytSbrya5OzVt5IOo4WGx5hFqenInOMY9Wca57ywhlG9pDYJ9mC3IKDWdqq/BxKe
nZ4NoUn8ywvyAOPMUhB6F9fL06D8RKs9MxOW72o8/MaZ9oB9o40LFqPeleasmTNEQo20JKVbXkxG
MB02JXKCg2ObuMQ6/TKDPo7PmlwWHITXqE2/tBj9IB52pWfw2mtqFh7gaYz2nvSdbY3/lh7I/KAO
ZLqtVKMwiHcy5Z/vDRRSS0We/HUdRN6kh3mF1QPC1KdHkSZd22qbHv0WKgCEGJyt4G86NE2Sg99H
YZvrwZPHvDDVzFV+ZTX2gN8H/il6gpd0siRLXBlauYcQ/FruSXfea/eofOF+YFYC/wFITjaUrfmP
iSL1XHv4hG9udi+mlvpvLc9BU5ysr02lzZ3/iY4bwgk1Am6jmLMPkg3ryAzLpWfff3gW9yRU6dU6
eoxzrdQ20METaeCTgC4BFoEqhu2ZKn79VnRpBGL9IiUKKdiPNx2RqzLGK+1wO4/wYcahIK0c4RLd
lgumNgxdbMX7Kqu9D+qdzCWz0sNtdZeF21kZ5CQo/59wK0UlaGL3ow/0DPx+M0gkoMI/YoKL4Ely
6O4wGQJdjgqySAW2k8kRL4MEC+pxQus1jD7x/GcmstZlbLtFiZd7pySwmbNKutCyL0E4/oAObJH4
745ggH3sczlsC/0XDfmBIW2n8x4NHdhGaTXGKtEJVEkUUnLH7wch6KY8vDcooNEC6OUo9eL8o5VR
7WB7hHNgnW3barf4TydK/vjX7RS9Upn8wMIkBOC2Xz/idY65vGciveUVMSt8pVyVdVjJX54idMac
ptKJSKcb3HC4MS2I9Q+YL3luALxJoTDqVTPMUuldDSv48w8qFRwYWMtZNrK1hsp6xtKtQxv4nWVM
aPrZ6cca5dshElskRiITQx8KOowbuIlvlQpaUk/U32BMUek0E6o2J9kjWmHO8LT2rm9NCU4yspF0
t7FfpYd8oMUUk1Y7AWMgZ6638Sm7edPYkWEtD5QAfid35G3jNjgJ5pcCONfYzdOEimrpKuDa4KTm
R4vhz+B12QLBUVM/iQ6tG+WPKCme133tp0c/ue+3q/0eNc73rXGoPH05mDCMix68/XwoQ3KC+Bje
hH4EtniLcQE/viO2Xdt4B3+WdWWGSCMu2lOPeSOqUDI9PZnkcLGT31FcnTLEAGxnZcJZ816kIZ+Y
Ksm5K+JVxQ0P+QBdwIh8TkSW84cAFjJQs0iM2oZ4jy75syouUzahnz7f/KJowKuwU97DV4ah8T8T
fFD+dv+6Csl92+qSwzYRy5K+fMRwRV+vByun9/7aHtis8AWdkqlsNnu17l4qXAyD8Oc8Pb6iWhru
7LdTUdwVFmbYzxJ1YP0rhecQHeYBz/yBbn4MiGBmwKk7QjXzRB/4ntMvFa5KU8LxPfkSU4xAf2Jr
hZ39aa3JNAY6PYL2XWwarXmVw8ihGpAwzs4Fzt6cpcLwUJTRjhh1ytqqf8ViRMdsiMfDTmMAy3Qt
1vl7jIj1dyhjlApKMgmRbBlVg7M2moXChACrFIKDSHk0vN3TDM+X0vPA6wD2XYSDVfheoCXQN0TK
M+94c+e7VteUvs4ysbonWqkahpAQJNHs4NbgcvHCPxOH71EruyJcY2LrKvt8YD3QoKPLa0Lh1xFF
y6dJIR4h4v4lBJRsBwmyxoCJpnsSAJnOmcaBgnZt+eLtnjfuiv5enmSuwzpJ6K9/bSkQKW2GcKR5
9G/iInKFU//Mnbl5uRVP8AoEoLyOLIDRU+Z2Baz1SVr8K7/FL703+pcgBPyLza/C/loAIr379HWI
QMuMoepaIZohDzuHBPJ5GRswiMXvKaYOsEf3na9xjohTCNRRUtl3ESweCtNZkyexNSNyGGa9XizI
vkVJX6usm8OyCG9BhUbohZM38wXTgb0V6xk7WZGtFnwzzYRJLwNkr360porRnpRg58jHTaZYZfcI
7IYgqQx7rPdSLDfaikgLl50GL0bm5vGZDtc4OE91peXEWAzTXKWwVoCjT1fEzrKGmYP+E6FiNqRk
+ubK1KVOZCMXBFjw0KwI3EUU16vYToWCLFKRNa9P+biqThQawaw25W5iaux3/Zk1lcpvDfx36KOF
9fONpYGc4o9vXeewARGCGvbbDG4tHi0cDfLnfqErWQb27SZZOlT7j9qW0rcTy4+D0qbO5NWC26oI
8v3ANmBUR2gIkcC8xvSSEbGQPWX3u4mTFQi5R/xYzMB8Dc25wGArs8lMonhiapbwrZMpTHvWxFAF
K7shfGwU3Udi4I11q+KI5V+OpngZ18xGF8sM7L16Sek3MBeVP9GBJIjfZ59UMkKckFe7HQc25a/x
rQUYPWC/JxFVMebyxcWRGd9Wj8Lsdqcwz7mFVOF+6Igczfg4Vfklq3AAlGxC7unnQzgxvNaJ0ky2
Yu7xjbRp3Z8DNfSLKje2mkeEqrRE2YYo23IBg6L9Yq4yeDR0MKubKE86dCg98RmBvloREgwtUWAC
KrqCHd0XpVTH8hpI/Xcz1pIv5V/FtX5KbTEHH9iEG+WlTTTJGK7ExmSXGmSJKRf3l45eRaohK8r+
He0oXLaTJ1IZXP5O+PB5FASMTs6VvKhtoP9C8ylxxu2qKzB3JMiQ7OiUzbESSaMmE8/5K4LpPHbs
iO5AqvFwRTL6vajJ/EYtMy8Amsf4q7OKq8kA5j+pG+5ntVmiIROF5T7eoZk+0rUo4cyEqBYNDj79
2EdJIDFJevvgQSoc107Avwt4ntVqINdT4EZnSq8+ut7bEpFchZjMb5Q677Zt24r0hyVM0GtSO5pW
ExQBaDva/PS2IKdN/Y0wad5Rfk6iRRpoKXci/l4sitBI65ktaCI3yyNgBDKkL3Qy4Unl1V+K2ZeI
J8VnfGzhM6o1ojGAkKkCinIe0UtmLujfnX4QImENxYDqSAwlMN93zSDfZEKOoNhEtDhgrUEP9bHI
Nwl9U3/L8mRFFKjWy+mnsnk9Kj7oyw1laTota4cm/N0VAsP7FXO8XBPMiW/CkDymvosILFyoHQMQ
7VNozJxPEFkDvfj8frmEFiJNAYAZ8ULvt4IzIBPvYdYsUEolPKspMOPILRUHHczehPV71kP4nqee
O3KR23VMN7lI9Q81Gs1ItFXmtcBM/RzAdS9gGJdAcd2AvmSUmG3Uydg/P/Aw3Rqs5eqhlQ89QBov
Lqd1FCkjoQpNsSk0ankc5hYvgR3Kvbzy8Kh64i8rTQc7jQdNhYeOI1YMCh8w2c9FvNdaxkxSTTnr
quyG9jx9NxHw+RUVqUpxHMvPKFVwIkHQyXQSmvSmalVGHGvyTh9lVnPmqZj7GNkarlwUtIVocA2P
0VI5CXYeuM3HE6BEtaxSnpZLGq3ZUur7Xm19aSRVR6Rpd9+mQDV2ByZK1RBFrrOhBup1xEVTsAbL
DLOhExXns2yB2gexIJOEbpXGv1GEiOysHTy7fXpQPL9jHDk3L+VuUQA4Sy/pbkhIhcsRXNcwn0TF
eW088AfrqxHvJBhG48LZ9NXpyAsNoP5nRzXzzBjV84cGurx2M1oNvosKkUdWhWI1uusOT9G2pjXt
KxCNiur9S3hfjYWBtq5b0jXuud0aJ0hTzks1WbXGgjtfZw51QtPW1J0GukMwOnUeou4KT0+6M7Lf
YlJ4WhA+Gn8q1lZDjcDm4PLkSm534U2xC4+JRP0sUa3Jl1MVZjvHTLjFUfTf65ISfz+d28++j4Aq
lveE4J6tso7vsSzbycD/2Vfkl+GGIfuRE0r7vq9cMlp13cynH1tsCba+ryt2aY2kIU60Sr9OXcf/
ASwZDo66QxV5fYVMRYc2m8SlSDCLREYKTTZjy3x4r9dZ6RwLdbYZl/mqQM6jwUxVnkzMzf7PLmiK
TMF82bPfKCW/CBUBa9Of83hzmlUtESz4ohJ9g36VRU/IwIwH31Bx08EJU7cTGXCkbI2UEiR8X/V2
sZILekOPvBijqu7VuicV9M7+FNBW5gboJLpraMdjuoTNLmqnbIyp0uk5VmmBIzqvxKAowqpgtUWT
1L/SDwMF1JEa5lySv5l5l+/B0eYcRv/lX+zBGgrq+spjbJyoAIKj3le06nhVnq34tG3qh4TAKYqy
NqQjo0x7DPLxgWqgVVh2Ez7+JRXys7FfzK5cTPzx7g9Q5boY+DIbP/bWxwQCqZR1SMxB9Qe1YzQA
oss9Lx7h1/AKn9YJGw+Oml6I4IFOcNHTkRUNkVMl8Rq6xv43a3WlRUWthF69NYemYqMD6yv3pubg
x6zcE/+k+0tpKKqE9lyWMWb4c1f1qkrjl59jZO2HjhIsK5wocxDLSnVacA+mDluK/bTTczYt2gJw
zximiptRkLMBDA826+suoFsU6i9rtdkxBXSmA8PHKXylmWQi4jnxnrO8gevXaIVR5RSjy/yxmc+e
tV3wRUeFtrZuLU4K6LmxIftIdugxZa0BOtt47jwC64tBAiHFqZ84MOB5mAtsUm4BIOeJ5787Qjg+
EP+NtK+8FxauzIPb2hSgSdPtBHUsiHkLgQyBXRvzDop56Hnj3Mu00xekornOSgjHAXpA2e3or7DR
u5WUdB8LYdahsrbfHFHvoKgYwSKnYTZh/O9FG32jNs9iBnmZz8alV6z1PARbme7SI6fl2ZzLAjre
SqMpLEYcm21EvXtSgmt6GLKZpeKYN3cXieL43iS5NXiYZ+3RmSpayfJRc2PSJB7uQn/zyxYDkkI9
Ec9SxWmrY84v47+0vHVYl+1pPiUi7QmS3YPptpPCIrI4lpV/GNVNZXcnKLZ1uCPOb6oOQpoe9znE
on3GkoOkn+lwI5suI6kjL9QDJCjS/oePuKP9mYbe6svJsjRehz67b3PT6e65EHFTagS+8+zJYVEY
SqF0OI4/wRlhgbO+vsE+HT8a6y6Td65ZLDWr5CYzrMvUij1lD7fxWscKuVgDx1br0tZiQYEvks/z
m/Hr1nVmZHN987+iv+Sv/kitFojx/VGURLM0saH5/cGaFUyOBvXOiB1np3nvY9j8GLbRu+Pah5eS
uQT7ybO8JKK7jaLPoflaD6JVoPB8iiyA0p9Mh4tLB2bJ8OjHL8yjKDW414J5FyI1OpoIGw5BgeE2
wBwrTHcWYJLUEZhlibjjaj/11D4RZE6iuOyGtV1+UVhg+IBisdW4dEXXT96ZPQsGJFBGBkn/z4pP
z2FK4XFVNuvt3/EyAv04lFH+hsIfHlBg8SiQzqWtAyJ4qLYbMIL1Rq0/phQGJYknjPUp41gUXvA7
1MhPeBJkWEbS0wnZ60We50mTJgZc+p7AMq84y7Lw7CR1NZJp8goBTtS8mmICKbPUimF20Of+GV0Z
BkX206DrQk1QLSuAnONf0jJUscALtR6okuZJsVrGkQAAC3ZkJRpmdMrVqZVYJWbWAixnbiNsbdoQ
fNx+K/X0zePeRLnF7ijGc4m/w9RirxQ0lCy6RCFq0lGqcRqi1O7W+X8QqlozlftJcXzV90d3v8q0
zxW9QmIdGToKx0FOhEyfP3VPGntflURi+NTpiplUGGnLMtUAO15tZTN70ihK/tgLSYJg18lJKcgC
WGT/fA2dEYGtw4h1u1hwopELC6bfRdNQUJeuisHn3vhF0QbVtJIJ68ouAmyD2AEIodcxTg5U5d/c
E+xRaFbSSolGNlGY8gvU0KX9+SOZBH3jVCSyjITJHX8r5gr4Eb7RcOVlFxlc0hJYLsqdC1zxIyeQ
WG4S4SD7pu9pDvJn1mBfwTSuC5NXPW95NoCdGC3BafOhtBf6ItMm+A3k5qrkjNmCkvUjYTfmpmjZ
R6AE6jBHtDsLl11t3JPoOXWFezS/3bNOq/ygb+Pcmyhb6pK8KI/jH3KvQvUWt0y9yFiV/pz4OEWI
ghx77Q0XN16COQp6vk0Qv/dPlQTTlimW6EUORpr6BVWtX6TEqtZdp+dRXk3O9SIy7yNaaK0Go47I
vYndGSwNe0elmF1W1SGvhym43QvXTQ9tPXCOXrFv+J+MSMgACyZ018RLbUsAVd/635YPQkkhR2yT
GiiVAaKD0eVGLVbps1gGIz40zi+7e/z3t8AfUUeXw9EvsABW6MYamY6Zjx2wHzUki2sI0X1nkpm1
yjs4Ztflp9STjQjVBRDGgex15OI2Ilet2/qF0kWUwCmCl59uLiYWzNt0qeOkZEP2H8bN5VJTJ6Mh
V7r4QPKk6YfzdRcNYqB4cNSgYu3LrwatpRNc/AHK4Mxtdlpnm0zDiQmFOfYziB/4ULHgxyGhyKgt
fpPF6/JrPRjudcdS52adXcb5FdNicf42JeIlG7WBLZExA0HMJzn6QMzT41bv6fVyKU8xelGlKlhy
3emtL33uekb6ZgqtruK8dI3Zr/aKSbg+JS8S/wTIIGpEXlJznCvLc+RBvjQK/FZrj54feKgbvlZZ
izfoHJg7Hw9VuXOnXzIWj4IeBm24jwCMmmF19N53KpGR4swDw0IuGLv3pewhikSUYv38EZaUeRXr
VB/89PP7VFbOO8193P9UaOzTyYZ3QpPPhLRJhoy16Mc4+S0BqdYiEK/eTZ2oP2wh4Ir15m0g1nfp
YHWKolYPdIiYlNjcqOdZJyNlJF0wTErje+F63zuqtC+J4qS+lX4CoPDmVONkACauzVGlBMal2VXM
lMl/UmLfmHO90c+Yb9JYMSCUQMOeEgc5iUG9jZOxqXMZ+8ckhJ8Voi/jgEN+D8LWv9BkRN90eLTl
ZkF0xbN20rQy9/jbucmVD2dURnOdp3vi8+lzEzgrT1lvpjJxXec8WqTKyrhjFB4T7LqVEhkSiRvQ
Qw9ApE0GEJq0K0sdav0iqzzRF/8w/5OZhZt0V2uWQD5Ia/CeTpoMSntAMDxwXG9TKZLdRuQBnA49
yfGslYbBKajOBTMEsiI164k6UFvKvPbptAe0W8A3TOgMDyMnIw8wMsD8l8xqCFgWnvjK1fyTtf+A
4A3id5hQl3Y2xCFfUWKpBDWa4nh2Vx0Wev0TnusCZ/Nz5zLcAH9mk4vZdVee1cs52xGM0sLUn93o
yvH+fiYS9sjAoClXdTtyG5Z5Aa63lFp6Bv+I2F4wQME/mrZjgT9QoF09Am1pBLkCGDazbGKB/eHM
YZ1zGpusRpuDs41YnIzPwXgnPMlUIJglwHIXHHJjOnNvkjv5HtjNA9MEWiFeHXV89UgUBWzqNwnc
f8HYQQLB9rg8RXNAztz9CcL5G+Q6bddAFv6nByt1l95WTn0QvrpBt8jEJXqZKZ5mlcKM0ST6pcSW
ie43CcyJQLB/GuZpebiNkI991fxg6X/F5fvMQIBJQ6VGykRDtqmkXfCSZRVRhwC5lb9uip/NM1ny
52b8MiaiVZf7KliXDk+E8D0In74ZRpZOLUcVv+xJq+hZ87WWaYQWgreqDS773lf8OcE/m+A8PClF
xsBXSWcUi1NeXtgm5Itdr3gcY+iQIuNSnnJRiJtbEz9RIAUQuh89PNmobHWlfzoXBl97fYXRPKxr
bxiPb78CyFT3dZ88UaoujdSSPTZDcYUnvWp4QHmsbI5maXAMa57eRSbISFQlGv0LwiSjJFoHZ812
Fi1zmG8GgQQZSHPdBeWEEPw5E0h0pDxxZ2CPV68LWWHO3bsU8vJJ6sMkg0/Cs6b3TSc33UQXtgAi
isT15EmVorTEClw/MijQv1f7DhRoxXGWHQdcOpNHgLpqjuxAhVKtM1f27DbwkmvvB31klqdJ7xUq
agp0TEFIiRo27VAd21/HdkqYtlvrymMNd5+QHAEntZTeXrm7OD43yvd3zXGVeNz47tDeGjFQ1zgU
XDUO1wsT1RZbAIqs1Uyb7e7JYEyf60tD4EI/2vkYfsV8yA21aFLAsl1oEbKZCuapZ1wioT5M0EW+
0iI6dw/mAtfhzjQHB12nRDmKgErJVLXyN0rWSlEZHMijIbPf1YdN2qhnwyozJalD86S02m7kFU9F
7gmZ/5pftLthROdQWbjZty08yb4UFDShuQZHbMoENFwjscyAI16cTzKfn7T3AYYLi8B+5Jv2ArqK
fcWpgvzGRTPuK+xhdgChz9mZnpIrTpIoPZ73ZWPuQdGlllfaZS1zhgW1z2ll2OLMwdZy+HtWJ85I
H4+J2BRBw67FX0ta/84jJYEJgZq5uQ6lJ55/uVDFK4DqD7cjsTZPTlUAIrz+7RdUO3tQZAFHW38K
I8n8o6bWTFfuuta7Yyf8mE/iTZOIiw14zuMMmZAM6RzFmjXOHkGHEbX1cgTFtlLrLRZTibhTuAm7
vjO3u+G0qdbLiTImCLUT1cNV5JWx4rK55FvtjeNH+i4aMdmS8Zlm9xgRCMqQ7QS8RksSRTbD5ql7
M5bOjADslIO2ZQhrx3Re09bzXvMg63h4YwD1LxBSwzQBVcQ4PFWNQuD1hPSaPTvHHTN7N+pQtjxz
pCwGdgmgSRNF7DbHugRE0Zw+UpFfJzEOSqoRwTNZHs5BET+OtCoq7VDOpWb21sepi2T4cd4CPkDK
OqC4pES4jz3WnMRvDM9nSAmVaR6djip6M7RkDhWs+/MYa+C0E3gpuHF+jIBP1VO/pz+2T2wo3E/Y
ef2N/XlJzIGiCoBtVKFV8d9aElyXNaVrTso+/AvxJT5jbU7vhXdV182sq87O1toIzeQh0Dxc1FZD
XmX78BFyzOluYmj1jDrAUSoPxik9nr8+X0rr7HHxoqvwxQkMTgR6Lot5hpDz/mJrNdZk8Mu8YzdI
Dc6sdCFTFrYUPSipoAfTPlxjaI29ULLCx8dj8PkyQW/tinZSit2m1UXb12dD+8YaCzJ7fvP0B3xK
+8NENmp54weqGRx2DFXebz7fFa1iHlleV5uhb+01bDpjl4Uk6a41Ffx6X/lUSFm8cLzVW1+gcHk2
+jPeaPXckkQDHtGPstHwrVJhe8fpGcy6CYxQA8X/kFCvht1jcLd0zqcTEpsjGIbjcU0cUbzZOLGK
zmHOasj3WhOYWWOFHHqvoxsjXmeFiywmJBJTB5ER7qDPOmXI06xudUrNeV3ecjBjOhSINPyNnHp4
XDSVhefAnqm0++5lqUNh5pszleYX2j+9LDeHi4fE9ydWhkVcJOgf5XrgiXcrBKbRgOur4Q7ZP0/7
lzTFMqJ7agym4LUT6MsvkXbYnD1NwX9Yc6elkU9HQNyn9FelfmE/S1hqbubVTpPBpjKsVUdcAjnd
Gwkxg6lCSZFHddMRrJaMIPox1FR2i0z2xL5EkODOTVouUYKpulj79QSnmpOrXKh/upMVsyg1rD8d
4Og+NVUEp1udt+qeCvlmue4h17M3GIs50x9Cb52YbaBN5PQpxGMSjHKKAlUDxT1aL9Hz9JALuHUy
4BNGgLhEQokwvuB6R1M+ico1doko1z8ZoHkyWvyu578C6VMleIh9FXOpF8Zisd+Z8ynEcOgS1heq
4qRvp0NR69F/+yj+fq0so/8Q34mRcOfM++RSedLu8DFYZkd8RwWTi+5hpuE2rhvLeSbxKT2o6aGc
MmIaWOJiIFAjXV76u/tL6FEbalYuQORB0LqCQnVlWEGrujCsst8ETxzPubY5Cyds8oxnN1TUVJwg
2kVGv/o/JWW2ElEE3aa8MBNrAhWrMl05jsUs55zmKhCKn3uhhE4XK6YMdLJ/qW1F67HjHYc27Yg+
6kXWYmj4IO9i72qXFWKIFKuO2os8cJMpkhUgZe06gIk9PHS+F80aVlgbin6RXw7ppFUrH89pUISd
unub4xgMPGR3l2QccyTaR4Uei1ZhF+ZEO32tZxv/eYNSlFkhoFnyBLjew+oS8NxmphXfsQlw55dJ
HC8xH7JxPOkj7FqUtYkfMUAQSIpq1ivfbewJkXsCZhHxLWeQ4jdvE1DzuWCxP7AYylZVeHMrfrRu
aJtGYWl7BUw8sTepjVyT+6WAZ50zk+Kav+5K4ypY3RKtR4U0HpWqyQjoDvZqPTLZIx6bSij+UkPX
WtF/KKPlGpMrNg0svgdFn9k71d43zQfwZ18raCFU7fvFoLNJCdtgH+jIpo0hNLICGf6miDwPi1tT
BpfnOigiRty272qufMm5C4Vjy9KogcXZZ6OPCe2ddAIggEkqWetOZW970ysJYDViKo+1h5jHPdCW
DjIhZ7ZuoOqLLIM9Hws0F4PNd2vPK7SnBMA8K+Q6ijkZmrRV80vAzO5x9O29YZHlyUx3a7Uayz7Y
R0fkl25VzThqppbsd73GooMu9XVNZK+jpEJh9StBl7qfdKH6KUb/mu4n9uNhtw+YJCGinPmwa1b1
HC8uDrvebdzvPPvtebRO6XNXEW77H6ZDAS/6ImLbwQMbPvSuncThI/TNfkvuWvWLf77Nf48eZ2A6
gY7bnRVFJA23WiUTSz3eNvAsFY15yF331iU/lQ3g4xcDRktDm+1AanmnPdtETu/d2txXqMW7IGQW
E+SVWsqhjPNkZUFYha4xsJw6ZBvbtkJ6VezAZvM8w+2nbR0U5kE1WgCa8yQSBamn9o33kvlLe8Lx
Fszgvm5BXXJSgBW+WtK+Ntbb8ibIYZZAR5zxut3pi84flGLROoS/YJOVZgQwdvVbB6mbCeDZd+ti
6AbedZIZjEbbqWOAvWBIJ4swIb8wBHlNWwq3zv+SY+bpa7C/nwxveL4Xt8vZQIbizgNrRth5AdQ9
pieNjdyFZyCvMcCVSIMXlK/qsJRBObpmH7zCkw0RzPVPj9da3QWpjfDqgaYFejX666xlUwj649NA
QnB35PA6tmlE6HtpUb556XHHAecRyQ0EqnH1cQYGW/cKULDObKv8z6Ghz3hSxusyqir6CA6P9NnG
/3vbWTZgz3RiFUETvXDbC999BBDgkPn2xPLnoz/NwQbs7w4NJ5SXnmH9nRqJ80exGJfXOFQd1kwV
XXziVM47QGRvWmFFWzq8vHuDsp4ZeFoL+JvIL06rkmzJWxwIMmQf+RSEpqqFg3r4ExfpuFGRYsjy
+w43Q1u1xnSfGlz3Qd9eUb/r+J4NgCKMmGfEnuK9VAT8BFjGIZyFmXwYiUKtkDHfu1AH4+CQ4VHR
q9N7LbAQfQTNfvja8YcvI+ui0XzjSH7M8/3LMlXo3Ox9oQBbrQSBkYOrMh4CxArP40R7/yFcTupU
ddCz/J6GPr25RXTbvA45GwC7emXsRl3ScVWwnXRRXsay6H2wqay0W7MpE/oabvco3ew1eqmII3+6
laInbkBaLmFVuWrn7bs/ao5bZP1jP4pPfB6FWVOSA9trpguQujKgznyGB5FX6iaJTPdBk2aqlo2/
UKoWtIYBYlSrOTKTTTtBldoI2EnlZ+Zb1wPA2Hm8elwpLWD8AomKoO33MZWphBiAtPtpiyyZtUx5
SmH6veaCcgc8XYtKv53eRhTIe619KXckxtvpZsj1Bcj62tMt9uSqXz0t5rojQ868hP9bTZddR353
7hmVG8WY+t+ZmOp2/tZH2iYC+wYUojRTkrPF9XYHGDLcKqLbRvncdlEPyDULeU6yK31L1CfYnPCz
dWAau5fjLPwZifJAzZJNyykOgVj4mzyTvzyPik1OmuwQfjgG19SEGogXm8giFVOBYGWkSncETaMv
n6GvMhIAXcdfknwxu9q/74EX/cZ0LdLnfsTgVLHspkL9hkCrEuL2cYQT6J+WwCESwxzsab0E+qQx
tdoE7ie0fWj1xQX2zVBK8MUBDIv3CSV37uuZyUcknE5HaCLVYCOp9L03JN3+PKY9U0ixTn8eiE86
Mmz0mfL4oMNgyv+UPLR/LZqszX+FsMpB6QFjh9V8D73KdQi2awR1DGLyDUzWRsioFnvfWILwlGbg
USuVx76XYRx3dZpUvE/jxqiNE1lFhfQFehYOTNBXbZA6QknM589nhXw9euIezGNUTpwKY9056iY5
RorDSDMfWSr+tKwNVjzgQ8TdiWdoRTFC4qtugjkgbqQ4HF448h8huL/2eniOUYZ5Xv2DJQt2HNuB
V0u85Wc9Tc9M9i2LldG+Sv5ADSXMU5Y0jh2p0aK9ZpoKdZvREF4bBVaxgmEm5eRqo13Z+HzsMM12
glQ4GUVr76gCOy6aeGZQ9H9oR66WBYlfhrVB9z97XlHEM/B24ZPn2JRXicD93h/c1oCUYzoVKIcp
qzLEtcyehv9UxCCJSaIyWz9hjwB0Z4EuqWnB92aTO6ezW2SmmJZFb/FzvMDvP8Wx1uvhspbzrg4s
eolBMrQZtG/W2LZ4oG7Wrk7PPSj+QO7HmBG5M9LlTTY8G8Z5QGE5UHdboZJHoC020eBGdv2+EPjj
hj3PBOb8fS1n1BBK0KNlUYkgRBa3+BYD73b31ihGB0udS8pHMCv1usqwH9zScPZpz8CayOGEIYDK
eDvtwA7Rkf4rpoMFUtrBp6befHusEkznF/9JK9IMKVywg2aoPrHVjEn+/2P/1+0jR1Ejz1VD1VL0
x3khY6EOJGyFIVbFlq91zwIcT7V40S9ZHhxZXkdi2xkFv/1oMWzsIG+QdN9tE72FAMtiEzOA1E7m
q4Q8U4I/E2i2p4pG/QG5PrzLbK2qKODwe8fuqYuoGZQL22wUDcQjtrdaItmKzdjON8WmzygkRvaf
7jcs+k7UsJY/q6ckbdAML5l6u29Zpt9lUweF4JaaW9k0v6hNFrLD/l9hK7tz4z996pRO7d0gQpGj
CwAey0E0cigHs8sD9PRgKjAOx35paUSlc9JkD7Yeh0IXqz7OPMLYlt1HA+2IbpWLke56HhVUPBfI
S8U+KQGLFNVbb8Go9Cj6lkJ58qmElEETgFF/Gsd9hkbB7CEi+uGNCYE7gb6mgO0gNjqgj/GEUu2D
Jz8VARw3cA0nS4cibT2imaFhxMDzh1xE1J9ZQwaqhUcEeTOI1GfkS8SJGLqyJB/06hyVi0r5kIE2
6wvul0OCuJqHdm4Hza0b6Jjg6mEf6U+YIC8eGiAS4WCNJcAXYmuHINaNOuirCVkZVgfdUsbSvxAG
tGZq+rAogakTR8H/u3M09igMi+nYxh6iSAOq5oz2mGccsKtnB/9foBIhQntkyWnvx+AJzTvnrJlR
VNOtufKiAk7lnj1Xj+GXjPTN5fHGHS4GPWuekHct2jicLEGHNd6ID0i+Fp1/mVJ5dpN4rC8bXud7
XUfAxNyw3cpRdijNbmH3x8iUfTlOcnOod/frhC7bsdcSeef9MxYFyOugJiJWZvUwbVWFrqIk8oOf
O8gHWpqH6t8DM0QmynhNBGU8AWL5V+Hnw6XTr4orHdIYAcyKeEMo65np5Qag0/P6m8DfzTqlB1ts
NSLrAyhW9z1LAbke/VSbi5a3Q0VkjHgwDd6s7hqbm1EMpTUUNSVp6oiCXRWXzq/qGPMATQnH0i2A
pN8dh9qtoLs6DyfoTdE+RY8BYWkty9XmE9lWk1IgNWzmBm4FPT7dq7PABvq4WaX1iRj4f7I7w8lO
O+bUrBteEwCSTH0hVb6lDEs21irmGAzgpadOVZBgIYwcXXbthjCVOY8liOXbl/rfG3Uvkpc8zU7o
EeyuZ+VC2fdc7VpFB7T8ym9L8fyAtT3PgqrG8+b43LsM3FFc4O7BsOScnCNndkKBpODgKIW8ldod
TGRGfJa8fpxhkrju8nTQrnzwnoyFCVirwKLYCO3L2f87gO3yIE51nMJFBtYcYPP6NknUxW6j3LG5
46NbChY1oyRu8npQldVnRkgGRrrkgbKIOZJSZaD49h2PFUhHjWu6B5Ak5FQE3LU50gkRGxOPGAEL
Ol5dqurg2DRqPmjA+YBgzNIjb4wEvsZFFOuXyjJSk7X5B0RJ/oXrLMPlcjg4twq0LMOIMLUIOQk9
prHzb7CNZA4PsBJUf7DkenRT5ofhBFRJuztpq4ZDzZyaJMclrBDeSqKJ9zi9qvtZ5rEQSLHB/Ksv
DRxL1nlIDLtG1vObyGLnNTVuWYdVFU8/Kl8NRxgybexu7fXPnt4Chyy7edPZQVB5h4gzffa4EIqU
MJNHCC/ZvkeralE6BjbxTxbF2euWnk55uJpfr4cS1btCCK5WyxrvYqHfMpck+4izNKTcFDEkp27d
e9eNt8AXzQqoecfNh36iAOYVsWfpclDjMLsGaFugIgtRI9/bZMtt6qhi52eFhgEwLe1OnqPWXJSD
9M23FvcFx1O1xt6JQaJ+66SawO+Fn3LCsr42SroccpzCOeSJfGp8ETDc2csEO2fNH0B1vByYzxuV
n1H+RPXbwNwmN7AyOPOp/EBp1J2OQpNwIik8tpuDlieBUWaS28YoDLRqZ81ywEvJFdmV5BYdOrzV
ObzX1dtm+XlL1DtKdG3jFbzvKMa0FGoj1uHXIFZ3dUj4TTWcJ1ie/7X7gS5DhBMguDswyZG1MYJC
kWJG439kHfwsL9woDR+KNbu3LxaLrWAkasFy5Yg6SWeL9UHBBFQPAZTPiUdc4LvpIjQXb/qANlIa
fHAextY2KB6EOgV60cqDdeLlBVt5PJIQfMBqvyHq0iE/Mn8Xj8IgIHmtmGb24rXhbEAP41b6nnGU
xqFQa5fvEyHG8+BGVrzHmjJWcRc5cxynmuYBZnAY2RXX2Y8wFSS4a4exmUiueFZK1Uo9lGI7/CYf
OQZCHR/oiHJiU+qRGs1E733husqZ32okPjouYrLPkNim7BvbzI4DByMU+CtRHg36RXuT0Ykt0R/S
4L1whgWfo0fP4vmwPC8IsykXlt2aA0ibWxOq94dq6okbi7+DpIeQuG7EolNqOcR+qBulLtopsnQV
mQuo6X46NFF66RPP6C07gBuw6p8KHRST+rYg/s8tMY1Hbd698TqAinTjcu9N2/aNcK0AgTNuzDtl
UA40elOXfpbkj5IonvFoduh+u2JF+9Z3rPljBJgNkeba9IiJYLGUs40pdXRRPx4eyyg18nbNV6dg
3iUKE6oIOuLMOmTvpNiGP09P7BxqiZ4RtPjHBJFt7CXGlibKsm/b70Mw70jTBlfQmJThrJndM6DO
25D+dK4Og5gzbQx0uSsiKo7nbb6FWSVPnphIymspGNbZkXUFz3t1gDiUxbSQHh99gFP2RZ0psIAH
bnALgyFx6JciPVyPg9cyBY8fzMVuMRaIEsfVZDdsfdsbkDZWu7WpT74hTBRVzaQVqtRB5oeOU+kP
chw6g/U3HLe2XWDwFFaDi0wc4y2OzR2npYIFNriBksZ1uND32i6PPtrvhASnV8Aut20tdajmAfyC
i1/d7ZL9qw1sNR7wl2OUAhf416ba7LKCt21ari/PpD9YzZlanZVkQ1oxysBmWoYmAP2WCII/8yxY
eZeMJHLa2BcyUfkoBntdeIAtlUQ9pwnhsjpXkpTkeYNB9PIFgmyu+RJmsVZZ60OPf4RRi2A+CXUJ
thwOtELpn/XA/4mcrgjVgkqJQKTIarTM1C14XwxVBdaWbfgDNiz3rGvnjApuE1fukiDenin0S70A
oKesUu4ErEPI4ix/4ekliYFuc5/7ap3Rmu+Q23L2f7LFfqk1fznSq8Zwb69pfL3z5NSKDWezQZUm
bv8UA28tGapIYa8q5rxmRZVIBasqHhCb9fqa88wLGWFz8RCIOyJhCrDEYK7yBrBcALIxGTZ5o1Gz
o/7J5f3oJt2zX87lwBQmfXl4DO/YvyRU+clxOAtsI3/QChkB1ESRXXRr+sSX3k4YryHaplTXNM/p
mnNPBE42rt9ENNg4ffufLR3HnNAMFnmeIXz/8re5EvU934J3gICgqmCOiiF6Fw1iBbbFM1O40Vc4
RV1VWE3eyvXXRnS5DAbmwrEHbr+1aT1tS+Ps67tXe1F+zm6sh095AZ/NKlMe5UNt1qYxK1c48gsc
knII8AFZQt0vh12iLBiCjhyTjbwoC9idRHMneMM1gy6rTUGq8aUGsO7cNDhS2L0dB9K3zNiUxrR3
Jd3FYBOsLFr3YvEHUvX084YLT42wZCGYW2uGA9hBEBgNDZW9J87+Ahhm4yT21J0llmhPfdeMuya3
2X2Id/YRAWtLaqq6drhjo4jckF5gUbVw4gqgVIxLI1pJjs/98ncHT6pg5BuQy0GxzylDLDs2RhJI
SeX1my3aATZZyq9uAUKpNvCbLBcDdYkQIV8p4bzJT+mdC72pBXBWrsFvg6OgcfQX3tCVKx9clh7C
E7KJ9Fhm7v7ICB//ZNzvExEJFOsP0jydAUnpXHERbE8G4VUWZ3sUVDHAG414DdTbzsgiv3HmQiRU
kv2xuleWZXBFKduESqeu6N4OmfUgAcmzJsnQ2R6bTbW3EP9AAMIGKYtktcpquSMoS+TJMS9quQhU
IgCkjjmPQQCvgDYLPMVtg0TBy9CoA76ijcSM25HFfvxzkQcjGbB68uffbF4SBkgG4vUlnVD72net
E9Ac2TbK/06CBMAsFndQYY3SnY360MUmESoSiZM3eL0Pg65cmC+XLsNRgwG5N7/A4yOmmIyYdD/5
pSanhm3natf+qSzK7FBLD+k0N5mksmArtNvvHiKSjUqseNN0xFxRGdMgCidXg46qHWlh1TdzbL0Z
XE6IYNCxqIpYfzcVnShgEyKLyYdDdyKhcmk9YyT1XR6Q3/Zw5jMuAGYwM5ZmzujANn7E0j6+2iu4
6MUG7F+/K1hw9Xzw/6zf01ISTNhdGZtVOO9ru2LbTmdRQI4bkCJ60sFXbf/f6YRAOO6MsZkQVt+u
nqMKORzkxuZywCQ1mJbbipxzzs4KvKdlDt4vcg3LWgDHzHlR2OeuGzye8nNADOT3sy2XgLBFD48A
fwrCvOJ98gOM9QtED0bbjMKOKLEtvMV34DKJNeUTr2HC3NGtyGKEm9AfAXrdA4NbI8LacFpNK6zz
p/Pa0tUzONwhTPMT4CfcKp3CepeIo8ABKEAdM4hA71jatoD/PrPAkTqNGGNemxio3PwReBy3cDxr
AlK+BJ5j8sPunmoVmrM3bKOhYtohixSq5eILRWMFLH1Cy6aZyAP9LhbAlF83SGF5c90jdxEap3hB
uHdliwALxz958zVNSbB3kfxsiKEhgrZ+HI64UiB/fAJPmxxo2O//sjqtd9PvhwrgSdxbr4frEwMn
gytrLmHrxRSRHmrcgpSWPTGeTjVZdP+YaPVInB2L41anO2s9bnOd3KZMj7lruobKXubyYTWJs7LC
FsLFFrK5KGd3hP9oBocBJeIC3vy/zUmpYYni9NGmJXr5p/+cZkPhTv8wt1dOokUV+zHe2lXU31X/
hIHZiir5sV6Ktap/p8FsG9T/sy9ER4vuKHv2N9dKjP1mycfb4FaknE8w7rUeffmN/BxB8hWc5v6F
gRhfD6GV+PmL6Vh/tuQvt029AAoJ1YhPDqq7j57cUI2X6jxMRxrSHsDjZg0hupeZTP3wcK5nNFc7
AvQazGLRG5M3HVmUgRcmL+L3UYJqDCnLz8rj0qQnyyI+N4WWIrzx5dG75UQkzEBh5TwMrigr/Hq1
gS6EEOFU8TtV9BR4oYzT4u8wt4oDt9K+qdZikf1aILU81jQdn4S/FjlV+GDcUwWXNaK3NUju9RQ6
7gGroKBVLptI3Mox1fpG1pULOPHJqsae7sPEFYSiB+qDiJVJwd9g2pIziRVaVmiXw/pzBVq/kPxK
E7APcj/CaOjdi3EJn3CFl1oSc4GyzoDYx9LccKx6MnwlLaqmiKYmC2IOI+qwYMm2JQLTELYusVyU
LwsuAiL9SHNQzE236A/fE1IA0vIo+DA2CdWMYxkMuNsVk+upQ1flb1MgFaO9LLI205qbcaa9D8HF
jsK72K7C9/76k+e/hqpOoijWtUKR73YyuDUhq9IdqVSSdyA8OjEDuv1+yCpj2osvz/z34/3AcCL3
HcaFQ68Fuya1RiW1pfdVmYYEWrSM38IhqRetCXJ7hfjZyWgdgjJkCsB+KJULrFMBX2qa/3AbFCxM
lUWHzQaZecWgaT8KWXu+EPc7gdgHQFMe5Kgo/NuK/YMjndQUA4qXQEMlAIuS0ztZmvbj04OmDlH2
xS2GmDT1e9LiiWV2HA43wjgRyMwlza1cROpEswgh1tZqjoGJwCzxLrDRSVWEbonRs/kPixTm89Q/
183b619LU41s2b5/AVcELnUzOTbot4AAOOnEu2qWt0BcgQZkgv1p4lURdoelMULwNdsQZ7kvUJ78
fJ9qtVATKHeMhaAGKjCzJxK3Gz4HmejHrWbuFfEmzvWReYYUDkR2C3IONu4eucObTbLiyCeTg3Zm
6vAygpQisdt2YHzlUqXvqTiSciMy3KFKUYvXF/lHRL2VVzKgv5V5s+kGnfAfT0y+2tlpQr6HqL++
AjPBqOoYOFkADWTM0tGWz0n53Pn7GNa83oI8skhvi6SfRQru4c1Bemwd2PbzPVsQsCNy8QnD6n87
bBDU7AkJBekMNbyh+CN4ze4UBlU2/VPxAEm/HR6MMOahetX68oohrv/g8eY/hWD9ZhzkZ9J3o70l
ADTWVlW1/o2gbXliobS0jfVxloxIx6npM5MnFcGfzet7AtIcdZhVOpX2hSSeFFUa33Ne496RdDx3
aDk1cVRBsfHSI7KEPsh0dVZFIsHbtRgK2KpkRQyCQqkUAQVJJs69gW5ePKKdPZ9oO/fKM8HkhMSF
nB5W9UiC8rR8MIoXAGlmxf9g1U03BzUzEr18+Wgwlv3HGhDwyton4Z7wpPMXGaUxEBGErlcY5yBG
YhlYbZVYRFIyKIcLBBRp5IBmdvXmK3wi9BrJ8/0NE1lB276VuEaKCdEn2OT58tdRzt3xDElUAhrY
ijj9qfG8F6vrVUQ55ucS0tCaVFkt7BSX1EtaDNKcq+02qQ2XXtN9JOFiPcu9XBXrJ38UghsaoaIW
0DuECRZ0K29tMO5A1DwOFj5FKmGni6YglxYuVHJwS2GcyjrEc/tznArcZwhMz55t1s6BP+0lr9ME
wN4rNWnkiaVaeqjlU7p+J3xd4Zs6CfmGXyu4JNRPZcVWrOAwsWrxNHhysJ/xIzcKfZkt6o9s7mn3
sQv16Kit0BBgDmEG3NdGZi+s9CBfeotwf4+Rqm8piUlRzLYkHm9mGbtvSM05qRixeP9VleDgPfyd
gUxvtMycFDZmmayZYESIRr9HZh/2mqOEmqkCcdPEpFTM7vHbpFZWUX5VQFG1hIog7GZ7UzTm6nQg
sT1ireBFwJtLYSeGdSKWBX4i9mEASL/EIk+9dDfHCpP2j4QkQeY9DMbzvEhFwOFHphN5VX63hzS7
7Z8t56Xkq2CRlpUqte9m+5knbZ0iYzO5w8MNgpBXJ+3B2VeCuKprtRl4M8S5OiUEflyzR6YlUF6K
u1c4vKFf6Cen4bfKtOyx5a1rpFTcjyay0m09IEFp1sNJG3x0/uGCHd8J9f5LKZGIFf9+VwgHEjpq
EbdQgi5ZERSC2dE78KkrsQbLcgYptW9KBrmNBuS6NoGDRsteQO5YYFdLlXaZQWbBDWrKhrV2UK8c
vApr+g9Ylbr6IGU4XuUUdq6WESmSQ8yRSuLlwE6eMzAa4ixLK4gDaeYXZKMBtpkbz3zDhy4dpIBa
HfbWn5Wmtil3UE1uzJsV0Hat/JBN2KWq2EPU/NJefFuyYu66tPiYinBW0pwAjdkgRg0GiAk2c/Vo
ShKH26JGZHuuiP0ohvBO7q3ywrH5qmHY90/RY/0W4Xsne6LAgsi3ns+3lnfM/HT9bVNvXJgsFIdG
Kf3sg8Gyw1+jQgtCTeXfQN+KI6AT4NEhVeF4eoCENkwrUdhJOGLf98sjw771vAtCfQOzPHwkAN3w
AJeUYfybx7kbj+TA1dx+ivILqhrnb9FEVvq545xMuP1oyyQUaqBCIE50bpyGkkoiuzUw6P0LkMFO
OfAm6lgsjpeGvCXLh7N1+3Cil/Idu4pPT9ruZilyJofcDEYoTb2RXozJC9a3Zob65Zf5tvFlb0Jl
OuoygPMa7weP+9h2Ydkn+6DyPB8aBCit+u5SVVPC/rgnB87LCGKG1vJ0tzlA+BjWdZv4BOLsryMO
knZPjQXgX5juTQACaxmGchYaTAclVco4QTJnrOkqb0t31TmcEk6LgUk9GvIUPlolD7g/IfwD2fm8
YaBQX3Np85tthsu702mhvGi0V6dhYNZNMRCbDj6vF3zyRu8dh+Br1zdluDmEt9hkoo0Vhs61hmIB
6OUHD+4OgWX0VvaLNlWZS9lNKjtFNHnNEQRNbMCRMfewz1OppM+tcgvwMADhbs+oc8MxIDOiFSep
zGjWToBhLhfbqusAThT8x01pUSO+aVRFQ66jN9tQgtdFFxO8BUwnVKehSloD9wN+t7qZtZDF/bRS
coBEOu8Ovx2i4yjvK6+rLJQs3DtL12FNqzmplCKtpxqB0iOs5rskwOGTQ5gWxjf1SXMT0zF0ZjPX
QQkGGMduCjGwXsvCVzMWm/kureRrgMYa7Sywm0Bkiq6P3HxibIzuUI9vh8FxA9MpAtj9D/hNe1Ok
3iuuaK3zsaUdpvCfLU4vFLXmoD3ThewW5vV8LLt9U9W9XNtNWmJoQoh7wTiYFExKRfz5Z+ihCvTg
vSUMf9fE7OPDiLtZHO0cRkys3yQA4LZwv3nTx1YHY+9WBY7H6LE0Pn4wzXhHaksaIHplP6sLGYQH
F52tFGnysVHgHFnOjrNGEnFqqJF7QCe243IdbTB6jGO9lpnTvDjbkWjoS7s8f/rOJQse/wgU591e
UaFDRE4Ggaf3cwZSG80NrYUvzNCN6lHrebyeuAuYSp+cqyJQ6hG4aKmE3fwGJrRN3xHa+LlpG4wr
YIXU3EztDlh/n7lLuypfEI6E3jAkObogHS2gR8DVS07327GP8OHL0XUvsTHZ0Mm7+DqOwqmh3gs3
VXDSs6W6OUBAHuUEhHNdYeL1Tk4XIrOckbeKHm9Ro9mgfrzTq6fwzx8m32AToVJmq7th2XBsopC/
M/28lm3x6CPG4+RPW+GoBgHDiLZ1l1lu8i0ycjBqHHuXFLd0rile+jePBUdXssrhB1ln88ryUJZW
tERtmt9Ifa/Oh4GB2SJquMLOhkdIR42ofyhb6TOpBV9AZTaWGrYNZo9Yzc3S2k1DgT5+bbq67YZa
m+/S7iRS881xFMCMqq52SdRyGfJS+BPFcjllYJUY9RC1MsLhvEq0kE7mVBuq5hADr+pVhuF77xm1
S3CS/yK0ya8x+94cWegsaA17hv3RCuXwNf70X04Eui1KvW3+6x/+qguyi3dDdUZfuLwDRJLh2fUL
nb/l16No20ujLgXZ5eeKgWMghUehXAB7+lba3D+C5WYYFmAYTJXAObHJuGV7WZhSmMTVMhG/wrys
dqfy1TfkeDXjvXwuC2cvZMQ80v0GXS7Hx7+aYzcySGV8QHAbc1jZ7JkCCu6cOZThzeL7lpqoFD2o
1CQAx9/p6poQZWWBuEtKKgRRxR+e+hV623cRegyNMbQWlY5cEhAT8jPi9Juq8PxPFFfYhvawrPRz
oeqdqXQsOKLKct5BLxwz4D3QpWhRpCZfGgCpEmSqFWrXBGjzZmL/jpSGtE4PoNXUgd/IEjALyQNl
S+q4WOSsypzf3BZ02dsuVMF4lOR9QjsagvUjo76XYyAjJOdfKmLZZHswXTOQ54eRbPXCyyI5DsGj
0d1KfyOAFkQRNpLnFRzILyy0ZPghcstzXih1dZunwEopfT0a0WzyBMBw4P7PBwL5efH8Fy+69LjG
EneFZb37hwVgw/xmhjhuaKRggQ3rBmRtrURy5WFeshhKrjrvrO9hp4eN7pG4+wyiKOdrUlaIT2n0
82+mFDeuuPk0JBqKbcpS9uXFkXm4DYfhA5nVcLBuWU5G5MzKF9YN4jm6n1p2QzmHI45Wcbcie6qH
a5E/EZJv/DW5NMQTwZ81Ev7/0LtcBGXXtm3MNBT8aDJ5auLprM4VkwRoZraCj+RpF90JY44g/sUD
0AaTLmR6geFDwTfvYGXse6OSjcmEZbXe52ixzkYCLeS0Y3TGQQcDyVMepu4Ye7S9iwwOHyx7VDDc
29a4Ex4aUu8fw4oSjcBK8CSyK4kSsTNSOZXhDH/e1wmH52M1GULcpr3bnXqsCiR1Ebkm5gJw3kQT
AwLMGw8pvLWNxzW9Z7vxAP1LIXAA2OMADiPNHE/qLIznVf0IGF4RE1Nuq8x1/vk2M6Xac4cAkU42
a00nhw8rsZ7A1CQO5LfUccjwirMdfChN5TDzzVPUjQfEZyIKPNo4K3gk/MdGCxlxJYLH6lbGRmmc
O+ovqmNPoCYyYzFU/t6KNclKy5UWwYRCRkcSK7r1zLT6wPPICw4QPmqceHPEVeecR/RZbqbPSspt
uYGAsTOZyg5c3vhD4IIFlMXyI+w1aom4Rm+evx6b3pzgnk7+y9sA+7iHkc0jftRvr4E8oERznuLK
TXp9343LRWAVDVMmD3cm6GQabBLeVTn2MNzWqPWxwN8rL7kMG0+cgQv5DQmEX7f4UKZkdpYZ9Cp9
pb7y2YteeX0M1zz2XOc5nBbYQMTyupFzQCZ/qU6OLPonMUk01oR7ZXmwR6CHqMreiY2ouPyOEF6x
NdWsyhj4JWLdwC5JSRBogUD3zAIwz4rSCbunPMhTe4bDd63CjEURZuISYL39OMJ5av6/eIvRwSyG
2yb5hlL5DGVwb2z0ssgABEbKgDRyjGrfMIRsjanEYr75yXcI9X9pjD06/OvWSnGKihbxggBDhinW
bjmdwp5te1hGLctIZBC1UF0UTHBNPpJ5FXEm+PO2y+2RN4ANwdopO8LbrRKtERt4Tmd20m2djvwv
dG61D2GYl0YFVST86NAu7gNNrgSwoXUMfdShJK7t6bK2SySlN3idjeTdNxpUlILOW0THJc22hN7l
hu31da8cHPYw94sdHplVgY8SbuFm8/cewwEDhB/O9Cj1f2Qc9BE08GCSSxqdqKLzMJU+pF8I/Ua4
xLdJwoDalOUD3ZOB/yYkGt3jTddTnnNtXQDNIOqi3//9xJ1D9rpnCLFlpW88pV/eeytUyyBpodpt
Jssijom+5LxJlpoDhMUg7WvhJXbYEegtT3WPLj+y/fGA74k98Zx96ZB1tXv1qbppT+Wc26bSnAG+
55XnfuxZCMhiNJcsu6reyfTJE8JFg9IxXj0JyEj4phCMzcpFQCTEPvRjNnkLpeUuiE+4qtY+xKri
O2JD9zZDp4cpgmzivjXuGwm/awuoST3ZWQxUe5GEEHJqLLmy+WIDq+tAUfJcqt7jVInC9wonBwZH
94ArYBpzTnauSbqSM0I8f1yGupwcZ4ZLSWlkq1i3owrYckdxyRC60iKlm+luMJso8GbkxoNxC/Uc
uyYfPhsbbpqxveWyhwTZ3fqCmdbB6TIJzlSbIb2x5e1waucpUDpngQL/7gm6IxZs6b9qag2HH3ck
/pGv9kI0hvedY4nsH0weFYuKJUYiQw9UNo3o4Ff37A5fPq5nEh0LHPcfO3tn5DkwKsbpLIg6ntNv
oWv2v84/6q2LQOIlOJ+TOjhSDWjsHpHquwJaX3Mf285MW/hYCWGNuxQzMxcs746LacAqW7MNjiox
kv27O+uuwkpFPVmrahg0W1RaaQWfPMw7VygcD/6FsLDL7rm2YzTkBYNW3hVWpKKMWp1uKzLsomeY
/xUB23KKS4oBx4Nlf0cSc45iqFfsbLiJ73JdcmEhAnba8vnexp5S2/qAseo70hM7VFOJ68ilF4Or
a4Fn/f0FM+PB9rpc23kw3F+YisFvzPp5aleuAi8CSDtC8JtdRGYN9eXeDkopLiOsXYzCBH230L6E
vxF0QgaNEFgZymKo7zSUwEc/nOUr0YrxDLW/gZEFJNkB8MmpHBURxWJSMTDNiXJpKlOzWuYpoKzw
y+izQ9vh58vH3ggWhVdhIAbwP/UT8T0BPghslRSH7HufGouvN4NcstdQeF4+0A/VmG8pwJq4ketS
wM+7IbWT5W6XHSpQ3OiyaRGYy4xoCz18EmWRNWXqjuBVaSrKC5gBYMA65APb7uOzd9h5P4GUi3TG
Dw1PUvI+CslTKehO4v0ywuCAW3xPVqom7LWn4lEAcWl8EtITQD10OZlMqGnxoK21ygzv+6AirqOH
WQ6aScD0H3Xxs3Ucl0SWvgfHHRSEPZOtc+ENc50cREPFjBx3N26+OycWT58ZxRAjFrAJAYKvvji/
jPFLBH9CUua8xMUMmjqAeGG6y+I5sHWw2MQDlLWmx9vi/JHySP9RujXQhjNg0JA2p59rh9FJVKZF
MQvxUsWgwmrgcJm0InNgfK6rNy3C8OZp5doiM62dra+ab4V9WiDDBKs2B8pVp4MC6smejTGXYNbZ
CetQtPu35bTSpg2/CtZKo6S68g/2Z6XMe+Dv+9BKprZ50SMSByRyc+sz82MeK2oXyQj6DJ03b/SA
jey9TqBuQjDs5ebcxsp6xv6Xl/BIFk8RSHe81ICQmMVYK1NLByTviX5XxGDZjotiZLaDU+i2ehuE
om8xxkEzpnSfjOuksBhfzzpgwL9bStfKgbLXLiR+TyRtTE14xzlumpQuOUYKXv+8vtwGFAL+cdyT
ua+4rwBpAtnSDDbcZhXV0JLaqaj9ew8BNQ5nwVW+YArZkPXQQdyVWhG0Rqm4cz6mUErvO+lQ0jdI
LR67ns3MJLCs/KMRMjjViYpzbwFZuby4NBNHbDduw2SlELyyuwI3M5NtCAF2AUGs4Rl5Z3mpP0MW
BziSCMS8hHFyXWeRI9PH5ak5GCxdqTplfH9785WrdiVNEqXeVWa4q0J5QdoeeRIBePYymV3jYyOz
fMDqdJAcnHs/GAMB9XxcV76xLAFVwIN0Fln9Ja97fMrTjj1s9XBclScc5/iVREt0hOOod3H09GgL
9r/nUfofOBxWqbI1dzXjCd2sxD7I6c0Q5o51/lLiQLcULAzcbXDfAi4L1zZribwdF6c3covPcq65
iP58cYIxp8GVOfnCuCtAEzcwSMD9U8iZKLUTXTQEUHqHLvqqod+ieHXknrAYeR+WZ7HfTTIi8Mgh
eYXCYLfUgT7TpnkbtCh0ViRODPRrGBpWHTaX2asMQUdYsuPPA+QfULlF1qFJNGIFTjqBoG5hSZxP
qPR12Tw7MNykt72GLzGlb1qGTx4iNbjb0B7ppU33SZf+0defrbv6gqO1heSOz+HdUpTwrMAAFvzQ
IbHt3QJ/gH4OZUSGKGy2N37vvVoK2FHscFrAy9Ry+b9YIP2sS4WRq3TSdRd3LsMh6WYBs856JtZE
CPQnO66l9ekMuiP3qX7wQUydMFrNOXvYqw5GyMqdSuwH5YDHS0JftLW8WqHtnxErhw/pzOeVquyO
8aHzQE/P8og+Wez+4HIfYbC3rWnU14oaTprnztV46CB66Y5ghhmTGKlpVRPOIy9cwUXJjT7U2b3N
TNoUApNULOw9R+RV2vtC7n093VO5IIo87NM+AAnMIHbUXLZkmlZHDj/WgbzajbCFcpvJjAn4986y
fCsM4YFmcyPw7F4idJE3q27t0Sfq0BoVD1GamDFI3uNFyVKRrWJPGZJGoMDRJOs2lIsu+5tRgn06
B/FfFtxD4mW0i/4ojiUIIpdKIes+KbbpYeo07yhHcPQTel5XSc/it+jZhdxpV0Hh9mxEX3mNdir2
7X3CLnLoSFvZtYN4doeNDLEp3xLeczPjcGovUmTRplu+M6CnEOF2d2LAGL2jwOxyqv+828qvA4ZK
KlhTHkUPdKPCIWK/axcmzKEP7woFqhtfeJv4+qnba4TMUg2ZbKOGMLL34k7FtKk2IQDYV7bxtFoo
tExwZXDZR5ilZnM+lH7MjOSpwfiqr4dmb0EmO9PzMBXjpntnr4tr05AK5UUotZRdY6Ld2bSJizhZ
P6xq6HOsDk+uAjoImDv6jsblT3TJEjUosSzArjTkmLzzatjIEo+xsGom8rpSD6djKhlOgupl8QN3
rADr1txTLEdZkxbzJzf6j3zdDQ4ZLplXfbqy3diRXFVJqP0BS0gIt1qeizk7bBJdOJga6stkTN6C
AybjpEiXNztPNUqPbb1mqnlQjDnUK6xS/sKLT9ynz4rOo6TR0xKyekVnufb7YN1fQJlNNt4FBDoS
+eg5aiF76ztDCDgrGveOYqPRoic9l7R6rmtrs9nCQ62HIxLsQCnAodF/hbmRnZO5o+gjlXN4eVVI
LWBBvx1AS2yoZOn1+6IsavX6XdYjsVj+6LVADK2h6mkHTJzYbp2MAz/b8+wfQ37XYZe0WQM/1lHM
8MDn1sdP/1C3JvWU0HZSAvFfvyt0lrZyCEWD0SMGYxEC2dPWupIKCOuPSjEmV1HJeLL+3uL+XZJQ
aZmvuX/17+QZDiCcY2DK3H51NuH5GYJ3P6QH5QTX2ndzuvkyYuTo+P0d+2m+aZ7+KVyunSxPF3fA
NBpeILZHRAVTzGMVXi/FSW3Df0xmA8d2XVMykMokJN0cOMXlGzSL8xTQGNvGY4307riMDAIwXVNd
ZDQMv5hi+As9dDhXjs8QvJcG7BbNwEW5/KsXWdeRXLoJSY7EszbeG3hK0EVNFzbzkoMP34idur04
Bwjp3QjCNemJL6OFdFm/HQqwy/fzaAhk2gAQs7qMzwzTS0j77nlZ/5aZX8RU28BIyhb+89Hcsb8q
FPpycYfNifPCKsd8o5YAb9buHMhJhPwMlevCJRUEPmn6Xd/mjQpmjh2BcNxUYPemmggNXDoXaQJ0
kNga6M2ncGO7OMku0PPbFdJ//Ue7sSFZds0eEuGzVoKdU7+7ATB2rCnED0Uh2fwTHUsAhKNFEYwk
Js31Rn8Sa9maFt1b9vZdJBiIOd/73e3iJWdU3DYkqJue+t7CYL+SfxzhqV/MOFMMsZ+b1p8Cnmqu
FJPdLNP+EiVa9qX8PajrdikygBLPoNREj1BhqBzzKA8HHoH7rsduQgj/JlYTCz5WyOzfmCLQ5AZ7
JbQnn7uHPRG5JTzRBgezqLG1kuUWy6f+6Bk7qiOUbxk52wKUv6Of2tb8PVECjxsSUkkb69wp8CTE
CQX1kz7+uQfVUF9GLkVGQxfSRcylNVHmwezS0VHRp5EPQfk1dabiXJ2KGAgUG5qgNrT80sgT8eQi
ffW/XdA5kBCvwF4S6W2Oee1N9olXRc737YLA9BWwRhvko15iYCEAqLvWoJWdxaE7MLaWMmveBGpm
auxKHaAKHxqlxUT9rnmpPMYLohrh4m6Wh2UiYXUARWjhP8Pw1XnB6k2n2nCBPLzbJDmhZ+1oi6UP
BlA1MTh0qsU2wDHViXmyfBOpHyAQuWr6Rp+njSoumBjF2kqBBdKAO0uxD40uyZOuZ+zAW/U6mn+R
rthGe/+8yGcet/gxnwXoKtaOWwNmQ9cVyYWrYvkIj30bANA6MzKvDYzsh8kDjGwIK5f62TOWQf63
Qb+N5BIUGK2o57xzb4oNiCHIuHTgCzwDwZQVZKxSJADWGaRDJYcaWzfbdALMyThBZ5wEBTsZ7VKK
u1wtcJx5E5hanenxqefURYMPkyargCTizpUwelczKxG7PBgNSs/8jG7Uvg3PeVsTb4ZjrP/vI0pa
cHssLEGIte/Q3k2O39ZrfNCrvjAGi6H9Xcjfmz7LnU+LhJIo6uY3H6mrJs0omHjClZVXEoP5o1xq
+qkWJXc2HzlkMqDOmR4hgzLsk7RN3oQuaHTxLIgtMs6NK0YH4W/cRuZywMyKb3tppdtQD78ZkaSP
dIXQKg7f3dP6wpJSeA9O1qRjnW1q2fbH1M7G5TW3T9yOPhKQxZnKZrpsUDdyDXGnk3dJwExxahYj
m53hWtAcEnGpDhF0uLsWAWT96uU2zPxZSn8n2f1ZF26aY9XjqUz0gyipHDIu+SCp6McAC72Yt6qf
KPLZRrXe94Q+XCSKnUCbKP10TCaRrYbqqTwj7VsgfwDwfhFzoCq+zii8mGiqJLG6/iPIWE0CueTd
L8IntAyc/8HK5/HvR5z2rM+Auez0haGwEfg0WflCUiv7jC9g5Ked3svqO9H+RPAMLagYlQN+V72p
8ZexZb0ThwSU7+rYesbO6u2b9rQa2g2tpzpXhLHJQXbEp2shIKLWLQC0AKBv5yqosUu4z3Hl0riM
RrLakFhLqVWBJY51lgs7Cwvfmd6Uu2XAvV8A1Is5AYYXAM8/F8n2DP8bjUY3RPINo73/aHafGeHL
zVhFGx6o30DaSz/xKEMxqOLLv8yUKHKH5H/eLslynKY1LrXWvUrjd31oAKe5OVdIwZkcisMzn+w+
PxKlksHhVUcmTsgLOQFTmXY2YRjfnowLm6NpWWMTs916WjxgeSyYHs4UIOOBPbjyZWI+ABmxv755
NVPxCjvj+1K6pLLSWzS7NjgoEraOXRj2z8D1mW2loIpUaskiGG+Cx51mcToNNLn/Y+3XW4SZ+WRZ
gCuvJMyveDmMxX/DDQtz71q4b7gcVEmWt+KHutQttCj6aSY5Ddp8rLLFAcD1yhGwcw3b/qVSLkL/
As06prDQSsgbrUjYQgjC+cW1mpSys12UBNG6c4rgDazHVuTOyjz1SNd3hul/3mUwooyYaJkjvCZl
WNqpxGUIy8VXMYWjozROByb+vMJXnQ1JFTKN855T75MMInLs+l+CQz0ABxhEv7tkbMiYHGib4bun
32Sf8L3p3F7dmMA61mSGuIS6Coq5OMlCXkDcOfQJQWXs11ZXznAklKH8NMjzF6Blrczgb/wHr8j6
ups77knmZP7xeP0PkOku/0Th82jZFLyyMrSgTHhs8iEqTzZChsLkIC8A0iFAcQ57sSdIRgR2nnqK
cWN2fI/s0PWKNxzxFTwwwsj9x9EZ8whmIg94hOheaVemaGl06lfxNmqsWCouH/Mhe1oZoNcI0x/j
rKAAHUypOi2prvaS7c0gtVhMJjlETI1p0rEMc2YhfJrqkg1j6cRr/N6317xMyEWWh2hgNtxnonSD
zfpbVfmsMJCBLKqC5jzqvU7mXCOeMQFORq0wIEaWHQOMA+4wOLtZXOlRbzg/YGRGnK7OrkNpsdQ+
dk8j1PUYetYtmc+NkEP/qN1badrNBpl3ObpEMQwFqZmY1Wp9Xh47NxS6IeWP/ITK8IzNkQ+OFlK1
S8tnA9uHpqyPSfNmPImptHfa18f2HF7bWGgLhBnkcJMZjOlas+FTayoa7kFLlQUbKnGfPKy87zxb
84Z5lE7Ix72F+zPsM2vzKAzDxDn7QT2oYsy7yFJmhgEZdYyYmZOSBDAcCLUvAu6LvtMYYIxDIPmu
pwxgDeh63rCZjbEzOVO3jw31Qpek4bQJwl/YJfrT0eYaK8tGpphYrcb6TNX/2z5KR7qYToLFa3C3
icC5Pn6vkUoIR8oK9C1BguM5spUbyeCxIeA4bPbgvIVTa29CxG9cwjcH0ClD6PVz8hbAPzbyzyMs
o1YRZp855ZSHSeXKft1Qw4fmwaM/IC+YP84s2jzf1GCl8QxoCxpg8f1NV9uHP/eJIHxBX1Y+oTyb
5kbe3N5hjwnhu3DadwcooZWTe//a1cdmLkJnmSa7TLAbTgma5/+P82pxvZG5L+hZ4K5iddJLQvO9
+wrgaBbBYut19CI8pfSjILPZT9Ovpr7ezyx7ue4k2tppvy5k1oKAzAjjSzKEguIMlJPkHCq4I0Gj
9AYVlV6BhTUIaXxdEUtAQHN3TRp4Eh/jEKVIU7yQzQ00Na1jUhGnFjBkH+E5CrFApBs0AR2r0uHB
XIWfDQk+85dSNYeZALDINWQ/wwKZIxw4KBduNqTNdo30HOEwQAEFkKYMBUWGMbprpYMzC0qo7O/G
ROdz34IOZq9dLpBjfjl/hCdVgfYsC8vjb31gR8iKMqlCVH/FsDuTi0gmLS63S/83zaCL1OZMJidl
yC0cTOLjdEDqcrNJdx7GpjhiA7MPNdxOJZwwvSRTWtV7Elxhb5KuE+wH8+QXhavcg86ri8U9U0zP
NWd5Z3EBA5kJ8Nck8skkDkMgNmBqCWjg84c+4qRNE+BdLxAMlwyF05FmffBQ8DotVXjoFEpz8o24
gcUivVN7qVraZOSJWBUlfjZUO1RnWPcLwB8iv+zYGn2CjrjluT/SJBFGWF8BQkI13LHrwwgQf663
Y94ua9sXLy+ZwG1W9xVoDlOmPGu/JfY6K7KzOTwVce01ZowuKB4H/TJ9Dxni6bpozXEUKnqUzslc
hj81gLS39lpaicx12gHHqdR5tvQEJDw5ldnW3QiBw1qGGoF8DCXB1oDXySpyFXo2FZL03a1SjXCX
gY10n/EeB4WB1Bf+vdk0A4Y7NzTvgkeE9MNWTXqW+lR6lqS1OwOUZguQcTNIpCu2jdw0f12SOvNx
ZcdO8ZLj7KHTaGyPApQ6j/3ZXBUG8NqJTrGRa9CMAZSAInwww7eqP94VGTpkcNBEvw+cq3ktSg29
cYO40j4pfFdFsoIE3C+u99yenS69rkCcGLGHeB4QRJA9WElvd9u49sVyf3Qr8JvTZ0A+sa3P5mL0
uLtz4oDlkbYUZp1snWbO4UFQ9B1ZTWwIlbzyc75h3splsFbuSABWkPHdHbzN2K5VVz/VMWLbacGd
Zns+bTsn3yiHdOVl5pAz/L1pI9CZwYHsathiBg5EBhLkH4UumdMR2e5+scUc+vjcau1trSTqSrH1
aPz+2KjudoQYKHWo58Z/zRkHteGf0ICHP+ROVfqLUtw7/v3Bii6K5T/kirjWgsvlGRVO7/lYrEVH
Zx+pEpXgXk7TE9T5JCGIqgHluQnPCcHHfLVcqtCj13c7ixm5YxmKvw1SxZ0lp350H/pC8BXxdduX
8ht1voom1xuFzSXkUb1HYPDzs7/6pW/z/jwAUfJGDrm1xv4tc1dXz53EQYhaemWLeV4iYf5yZSk/
pUFhbYJ/+LimWOFTV4byAGzviRMERj/YIdGfEhxi0znK4mEPhlsdXsH1BQr0HFVN3i/uzMc0SJN2
LOrse+uTFoZ7EhhRwAM3bY5l1lYBb33PxHPRp/yiDYokFePWMbRELjkuClq2BzD/UQUH3tHLkcia
yMw3YL/gcQl5sSXK9MWd3QIK3I3JXoanITcG+bedbpgRk6nqqnJxjbZf+MT1Se3r/aGBFO76Bjsf
nkWSMg6duG5R0/4DubMjmvF+wxomJnHj5ca1IqRaQnXhDv6KoxdGR+ZcZDJCT0Ako2zJat4Dotz2
oV1uOqydx5+XfYnCkj3DKDSlR7FWZyC0H8wXpPko1XJRBYFs08y1v9t6k0iZO9R0RNFCRB524iIw
0oAlb3GkTfch3IIT6bY22jRO9Ql700latRXMZlX0V2AXGnfAjC2VcIZKuMKv4FBxOm921AyTWQSG
WvPNm24etdC1OWzAoZQYb3hAheBCZ8I0DP3WMPZbvSEGOBs69dRqwpbwk+cNoOcrSIDD4bfSLsXY
+jdXo1eY7C7PO+sg4dNJ3MZi5M7iYgTr7swltJ5ZP6daDBVQjbFvYSi/YyAKnAWr9P2Bp+Qj8Xgt
JY01FZG6Q4flUtwY/3Zra5uM3TuU93qGBYcZXYc/IoAWFIXD2LSEqUoOAyg8fMjdaPjbGZ/r/Bpo
glQy3Q5Nq8NXK+cK9jzG3g4uxwS8GsX3jMqMlnDAu3SwKNdUyMiJep2ecspo8jnD9etqGrwfmGkm
4FEMP7YYbCOV76UT0E6+w2mc+w0DD0hP2UzAHRJ9nTsBoRfCR+gzOSpXzl52Wr++Ym53qJG2DVLM
KtIXMzrH3BS2JansNDP03+sdTGOFLXPOAR2Coccb/WlaVW6hQ4E4mdVml9EmQFokXD0mJRF021cd
4AdtprWE+k8DP1+e1CsYz4uo5XqfMra/dJJGmmA18Qw1MWNgCztFLVZz1a/HPj3J2L9VMa4OrHTH
Qncxumbj7hYzknr9H5p498Uhq/oRMWQ+XZGl/hG0NJIL1tkToCASiLourK6QjHJBVZaQCo7eDBPe
wcHDAZPwdFZd3KhPm1j9N/a2K5DIe1Ta/tnZ5BIytC50NzFKuqBYqDyfVDy6kjWrDDZCgABvZjf7
q/sGrAJ7D7p6JRtTj14dN5gbI9hMxs4QkzkKsbtdgMrv0k6Vnw1EL1Pdr69MkCr+XKRfBvQimym5
HGzL+b0kDP1XU8mCQaPZQ3vx1yH0bex4OOonkpVz2UNYmC48/dmcWYa6qL0E97rofLehi31D3UwB
1aObX17dd3TG8eL6zUTRRsuQ6+KGIgeC1uwLnmzKi3wsCzjdD0infPucbAFkveG6Wt0Cn5voaVTF
107DGjajHF5Hr998HDsn7WsbyYLIV9ZaoZaNNZ6QkG/mhmMrCEHOlpVNwaamYuT8wVjO3eG42xiG
+9NBrs+hxf5GzOvstUoPHHmKRRIryw66XzFFgoysahLfahynATvqGYOt/nddLZW4Q2YpxPRSInvE
mDi7E7BTl1JPAIIGFhSx0qjDYNtHt47rYKrv1jxJhVm01LiBYz9meRrcLhpsA/NpVquTe0p4fiul
B+W0E+/C19WzTv1taaTv5bm+gzk3w3X7vsjEBgaCYHfyZf3h9pXCJTF3qSflmuqpMWc01m7ZZviN
LhHITwG0tlOj+fx4oUCMveB2yk0lblngauLUNsV2i+mxySh+dD8OA7kLpZOssSY6T1EEgD6JftgZ
5j2ByMsybhZEFGrCUamSNYMF88DOwUE+zF45iHWt7EOyOkfatEAK8RZVymt0YjI2LPVdYaKe7BCt
CXcA4diXnddR/oB+pBWr3j17n5FO636GcvXj8mqMYbH5qFRnu66JOcnPMRXrDjwIJr3Brlz94Oyh
inzQXN+7VgwMeQ8YEXTJFFlaUFIn56kfiw5SZxbBbe1Hy4484tWFbggDuKchMYlpu8P9YFzW8s2k
euIEizCtJQVfTVz65xaQWPh0m40mHCs3WyD+BiwS+uEviovm5tuZTENYxEVBkB3ifS9b8LRl18ZA
mAXXn19yUtFOF0BweeNshYKKy5M8DGv1uyg2lyfWxSA1KwUQk/cny+u6pml0wjLwTaNpFFtOhnrx
WJtJS9Q1gjxjRtWqYdfSU6EjQshDvLpGT3+PjSAhwfhqRR06IxQnmbBxbTgBGujCGWvIDCZp75CK
uftZlgojz2YRdxtS0VhdwOUq87LfBSv1dOBBw92uIXmTs/LvOez/HCoUvjVV9ZhEOJlq/iK8FgOg
w0FhISsFD+riDErtO3FKnUQSECV9wP86cA83T2GHCjHT4oRerw1UUsnqZVYvreGYHxWGi9YDG1Jh
6zh2YPjbcuk1osHj8+Qjw4ABd0RIR9BP0XjyzEa9/Oh5HX0ux1diryAXUjlA3d3qmdyLXq5R2CEH
HiHoPvu/yjgSLmdNPfHpTvZXLH0r2o70DUs9PbBSk+1wOIN4pSfqmzYQP10cUfN+BOyWRFpAN4TS
6YF0dvqDUfqkGETJcxMP7dUk3tBSx+hqsuM9woWmFkp6DNpODc5RYuyIqZMdHppKLRCC0pH4ceD/
4QuLqSmuAebQee5u1R3wjIhHZMcl0FwtLKIX4RHSca3ICKwj8eFqINvIVOFQ8fyLPJ02Yk02v7db
qdPyhdyru5fsnyaao2nKJm+mmKlOuM4t4PD3Qf0mkbcX3KZuE3dMj9LHOKH705tilxTV0CHQUGAH
putNEZB4LMp0dUOfUiE+k2tOPrv2gQin+n9kcyFhUQ2+gTD3c0hLnjHUUwLOp0gYaxzokkRR3KtD
m8hT2wkqA667zHtdbDiTWKuF2Eav2wy8TfqpVY8jfB9Y8/dK0+bzu5jyYoYiEsoM16vIgMAibgp7
11eb+R0iiEPIKgDkiNPuKsmmm5xEQEhtL90VChKW31+AbuLpk7TvslYmKKlbyHQAACa23fPTYxlv
tAXWXL5UAbaAe7ppw6dMFQxG4Wg3MGHBk11K14mLjZ/Wk9wu1vQM1YRVkh+sZrAtMfHKdKx+c1tI
AZOGfht+OXnZlexkyhirbb8miw/ibyaSnxR6Qc+3opFCNe2aT2uodyPkTl10v+ee/FoTknXQQGrd
iuZsBJU3mBK8ECmI3quPUqz0fphQqMu82hPKDYt4jjVh2sxrJrYugMgFYhFixxIB6v9bd8KEvPTi
BqT0Sj7a+uUTYUgdL8xAoLlr6A0Tj2TtsIVyXxj3lR3uT6lOYgoWiJxvgm3i9Ztd1QGNbG6Mibkv
2hE4MDzer72MHPZhozf7LKneq7IyLu8oi0132StJgF2j+4CzEXqCMhOa2rurc5QBTswsd4hlYjE1
++K6rhKQMcmLZQg0pCmww+2o0YGsnMjuEDw3ulRhBto4HtYglPZQMJY+85ObqFIyiEDOWUt9uXS2
02V5LNpzgq1Xk24b0wUzzp+mp3akbmWB4oqoJGGyveb1SLHa29lO1v+NbHHGxTA3njrKwXxHuqHA
H3vywAQLVLfBrhJtZGxG7q7guQiIqryQKKrAsO3AWDNiDpa5/iLtdFQU1PT3lhG0HQwXd33bc7PY
LtIQlTGHD1TEdfpqHW8IGpZ7aHWhYz0OBSBHv6xW4AXWnNllcHifKI9p9xzFHLVSe6K13oQxlRmF
lomomafukTcZNhBqCcFbeXsANnPTJ8RySTa9EAI+aIBUUAC9yqCjd9jV6TGS7oI/LN+ifgTJnHF2
38U0jeZkSN0nP6j76KayG3xty2VqCbO+jTjVJzew7J1dmM122/Hur1klTQXnLBABOsTNxG3TuzX5
CaxSHcas/ljCeA0MXSlSmGzqBCupB1sWGNpukgribG8eo6W7w1Es+8BFdlO10uRroB/idbbshAeq
fQEhUrvuGsqqvx6uMQhe24Ns9EL8sAaorab3alOXUWS0YsyYo4S4D3pzig4DMDPh8+AKo6h98LLD
CWunloNV6BEsMWF1xywnsoKR8vVwLElvxAcwP4ymyLpiOYWhKLJ3e0YJbIkba5x5mk+oqXgqOOvz
OeAgTt5wwwpE5VHZEUj/0x9dNf8uwGZCg4yXyqZWamPQVrW+4b63LN/EY+d3pXU7L9OhwqEoLbcM
9W2aNfyj/hNr7zUvWDRcsw2SRhVBwgQanl4+41ROu64EjfomJIMamMLMTGfCZew7UW9wBbQ80xg/
8dyTo1YAvAvupuuc0Ejt/YF9iC3LZftnt/izaLwyoKAGOnZxrjRndJm0oytAdPKYdHpZk5aeS3h9
CO3XuRaPSYAHu8HYOkvjNlwoSrrbLkn6X5yF1ouwlqrxS5nBFuHgSiugJTpTI2ZbBUlOCgf6a+Jr
TvOcHmvMPViqZivKEucCsluc+uzCkp7sFqM65wy/7ZeW8mryZ5LTX8BDtlOxbe7J9WOtsjQiby4k
WnL0zT8OXhXzujj322y2fEQgYono7vULapE4LaO7Smnc+EOqjiKsTg2mpGGbYczjdSpx2Z+E69MO
6ouaJ0WMCqpamG3DbqnKUdqDIBF0oIIy7Mc4xzIlXWmU5MAjSlSCjhKqaI6EtbQb8CCRyg5KluXH
GQ8dy6KZr9nY6GB4uOczuDM1oQ06RovI8fufLjC3OoRvni69EBFVonTdGxbU5tRYT1jNCBD8FlX5
cv+WzyjmoKMFddiUETSZsJR+0csZwTFgjrZ1IlUUcs0knYSW5rgmJGoeWpBw3y+LsH74Y9yb2Tak
I1+9t5j6KQlGwAeoJpgkEvPH9FttDIkLzl2egKRewMbxh6Zk4iFZ24DlIiaFvm4s4gksDYoyCyK9
LysFZabasC0QGZJqnqJbyw5lzkMr7gB1xuZjWIbSCjA6GUEy+T7gL5A/L6ZbZPeckfbtGlQwFkhV
MZgEh4DUS4jzGEHOX7DNSyek6Iox/iIGTpwxlrPLqsNF9AnWHiUJldq1p/v/Bp4HC6Is6RttY7xZ
K4r9zfO2NQsC4ShWV0y/tHLcd/P/1AjU9qbFiw4Yrpygt1xJkULPiS3JcRn4uH4SO4LgMwyfuq4S
dGIiTMBiOXyyiXwy/DhR2GmxuA+J8Ng46WsJowHVxbcrO7uKMVLpsKsPXIZfms9ZzsmlFoPKxHgq
fXzzAefeWdPC8Az6VpdhGyLLflbdTNngpDBUY2lWN7vRXtLKNWLHOQ4nWh27JFlchN2bjy1DQKLZ
yspv/d/0dFuOQjQSUx4qfZNTsNfJjBFENUxez6nOcO6/lQ1o/AbfgshWI6LFmwHYCZ3X809ajJpr
47fBEpBMQphYs2oez5nIsXzx9tsFf0v+VtEOKn0SArZiQKRw5xiseoVicaa2LQMKnaykX1XiZ7Sw
amlq26TGTFf1xIPpiFFfCEiHReWm1REVLyfRht6EHMdupTf/VzhKyQr3dYFo0P4c2Cnzlz0yYlZg
0Cj+sjhVWh6IYVJs5fYuAlkFjefmsL6oyQWQGPTsFHQzGquOmtcLKjjemSj+xmmeNQjEm15SviEW
2mYURXFQoGMBgLfbI4Td3fn0/TeCc9Gjwb2HROo54HJ1jfofyiG9wO8EqmCQ+TSwz0iwEmg5XGga
ZivN573VFj06Fm40hOsdzPUwADnYpasyiR1W0eVABhc6z4wcwjNnEPwTgMLqBnv96vs77SxQl7+A
8ECXgSxI/GNY0KI83rTS/bB0+eOaHUfrC/T8nJBrK//9iovKmtjfVzFlF9bcJZ3T7UsM03SRuY51
nSGM90Jw1L4sWQB/hbNibvHtWeilKAEmmWaFgQn/wPKYvpu0C/72azouG7PyZESzZLhmEJrTPw7J
fK59Mvlc/HrD68ZrVCuaRPSz3elH707J2lXBdp/gXuJNQt6tc7WAB0PhpYY80aD7skR1WsEJ0mso
BO0KTPjL8EyRU+qOb+er53ZOFJGyXaKIwqLZ3LZeekew2TGj+CcIQc5EDMUJdKiclvOtpfvBIehz
AvwfenfrP415hiz+s3SAcY4E2nfXScUaVIlekA4U46a420fKAS9Hc6WRPpfbXqeMy5bKHEaPijui
/gJdJQn0zPACACrLgVRfXU+P/PpvVPoNc8fXb1jQCUenhCe4gsWDKUifcIA8y7t7r4Uq6pNmybSl
2p/O5Dvho70voFirXLdU1BrtQL5IgrhGT4HHTPLjroUowA+1aidkXKLVdiZ8aRPV1Gnw5hMJ4S8Y
Kax84g0GH01EvB1XlYPHDgri5Zg3WiDAT8aavdTIseU5dX1+Ao9BFrryE9pEWBaFvhfpOmRXOwps
k4GMRnRPawKPMoVjS4KqZT4+4dzlJXtmthZyLkeMv5HhbLCb8ejtPg+usMjohcMc3Q/VSMqp53N9
640xu8dh3M+aIaFqjpkQf6CdJcJ4uu2fQGB0T6H9bHgnRV+SA4fkfEBjR4gYY0res7Rz8pPnV5Sl
nhVTV82NPjjwGVGwhwNX5KkLeCndUEV7ibyvvmv8QmPSvgy654XbMjllYMGrtMPyrbrcur1gwL0h
waxt8vq9CJKUejTgTWL9UvgvT+4GCy8Y2naLbqnAKZkiwmqrb5f4AH8LhDX/5nmWcQxkPLr0iH/0
iVe74zJNe7J4pOVb9tQDFJu5nwj9VvwkmMdlyNaWuYu0YoddO7D8lg/MnznJ2tF3IaCmSlO48GlJ
8Aa0J9n0n3zbyAKSP0c5HPqpJ3j1EnZH5c36mDF+tF6BEpv9X7SWu9xfML+kCJ+BPXxBHLzHGYnY
qj6xwLj3kd6XAJIlYj6kh4DB30xaOCcSbx+vtl0aF22DhvNiT6Et9uJZdKNE822jmhggPJ7d2bFv
vRZxNnqs/3l2y4DPffmp+zdh+uUD0h2JHmbxTZVWiwwq5oBt+b0oZUZ1hcToutIpNgPsRX3emzwr
n1JLS4By3TdoAgMF6r2PZkJe/TVev2u+Ur2TAgGSiWj5pmEiO8qIARhKmPFmiw8bcEqdNrEZ5ed6
I+fkqERi6SqK9s0aj3HRzgwAmwjDQy/1LEQ+azI0W4o+UthaSnWssZlt9mvTwXGBZ18b+Choe0T9
eSdMyg9tZZ0YjAAx8v1BevX1/vTxdbNziGfAURn/ZKUrt1I9XaDuGJNX9zp/fHWb6hiZFRAkuIA+
k+uc4GKbahcex9vbT6MiC9KUP4my/N8Lewlr8HbM9HGVFeya3SSwThJxviK+RGbLPIoI8Ei2ukaC
Zo3nUNUBuQuq+SEllhzk29U7AKOdE+D9npERa93ajwDejRYsJ+Ez5ThS1VBCyIP4qE8AVeOjYhAk
gUcj3hF0KYGiEG/eYb3NPPg4Myg+zHk1GLMnHyo7jNzVD0sgPrxE14JxjBmwUdd0JDUvHWILKzMv
T/LQ+GDjzCLaWnoPjaVQs+icphdhAtUkbdNB/HiaLRhb/W4Dpo6nIe3XYkOCKkeCuOKXspvk+HdQ
RXTe6CwH0ObWdGeIKlDcBLdwFWa0SN+R0q0RWcJ7KeQjlzeuv0l4pFguZlmnR9EI5s8V0n7uhpXH
qDHK8M7d9MEnmUyyppwhHnfp+U7yf529wuxEf+74UbewXB9kjdi1R3YDuGvlrR/2qWSmvCjOctai
LW1ntNb8Tcpsb8iQb9Gu37e521OzBmtPlfCZ7JkBMWc483T7Rd2QbuuVacY7C5qAACenJWzlxWxg
JOfgSv061ZdX4Fm0mtu8ppdSsTRiJbVg3QsktCfRYmkYcfQ+xKqi017H/t5AB3Zes7k4yrlaI6v9
ZoU700Dj/SBox+YX+oOofNk4LKReXweYRo4G9WDCCOyJaPMuy7DDyZBmUWKfJWZJsB+btkT9ZonW
kVUq4orq5zxkaZz+IhFFvVNTrV3H2HQDCl09FaUaFKIZ5vFGsyMt09RkrNv+2YebCN5oOAPQXoGA
CxkmakuEpV2uE3S49wKc7e9gokbeLRRFafoAoKyj4jDASlL2Rg6dnXJIsLcCvfKr4vQwXGQsH709
gYjmrKxrSa/Tv0EhYiB0GumBcmYR9lgHVI4ush5NJPyRbJr6Tl6lgWHvNtL+yd+1sjuYOkDVXJ9N
N7AGLw7mldWhAv70u1Mcwmgy8GtfInsdrurT5e4zsw5KxD5bh2gFT0f9TGAuoWLwOPGR11mp0A30
3sxvhs5iH096Igmc+nPfX1NcM9YN/yKH7jm8wxfq5DRUeAbz7FbjB5krWSJFX4j+VrJqWp5GOrbx
nXjOIVH+rqYFVwVhGupRdaJM5M3gPp2DF+TuywraV98ZAseuITiBzWnrEESnqOgcty5b7+PKus93
bKRTGl3WGh8VRm/Y94VHtRVa1zy89qplYv4B2nZ74vP4LhYDG5Th87MNv/SQakNu4Ei0PkiME2O+
qzO/F6govO8u1DFFRwMYeXnDqxQ1xoZkmHGA8a36hEZ6+tHJ37vksZ25g9ILuJsWfi5wwEIX7JNP
PNqhma1MlHrKMz/rT6WXaQruuymynOvrt58XtKeCakkZzU4vlSL18fOwzrAm0HzUJN5HRWFtA6Si
P93DDpTmtgvLsb6iVhalsenA4A6Uw2gTHQdYiCdGcIpjcxIL2oOD5ERI/CAO3kLlGHJHfjxDKqQn
f6mnS36TCT0UrAZSfmCCDm/hCFlXXGZDljE/28o360S0nnSQOJ6WIaCP9+Vc0a5IYQ0VXcHMbcGD
F6LSf010x6qZ5hUEsYCGDu2x6PBAWBh6bSsNF2yXJxzbQNHSUzPyXg3FSdAUUoF1D0j9zeYJJzTK
OvwwJWeOJOD3L9C2FD3G5LvdZhazL/fiXZPqvW+RjfsL3vv6DTBBGENt+beOLmO4El9bDs9XELuH
hr+wKCxoQtN/LZYmOrmobNo10PnHwndLyeJ/vH0CS4IjYSepQoUn5j++6sqMrvl/u/YzoHpzz7zh
XYsJe72s2mfiri4wvzeTBK4e+h7zk35ZZeszvbcp5MBhQHYc8ObrY0ZPd70/kGxEaeCvVutVpdCa
qB8mwASobMj/jyfLuDHcNu6CyVuImsjjQH0yAnA3O3Rk2bCU1o9L/YLYQpq+rPEpel0tPvtdjayn
KgvXBLl3YRnZxIYkBX7RWj9+WR42hUmcQdTdem3fuGT0F1TPe0iAe0HxhhosnICaRl9Sk92I02Vh
SzC823eFEJiFKPvAF3+oapdvcgkf1063g0g3vOJ89UNKWpJAd5aoJX5p6/Fib8jFhv/fjzec37Uf
pyNJpGjTJMF5MVwv3rVATcTu/j8T45GWEpTLsFFzoynK6dIcJ1EmTPzDui8osAnnMzY8dG/Yjv4j
wtTGNS0luAsDcd3ItQizptntOHUGPHw/87rdp6TZ/TnuxzFtstDyUDrTh5qAtXj1BlsT8dtevYQC
1Bs31dmyJhIDm+pKwbvXtMj3A+SaGKiDGMTndRN1ftZima3adt19UETC81otyORdBjgMpYmzW9H0
bQSRbCEB0GvAoOECcBoXsgXIg/tuSxNpLgidYQFErebGydDJZxQZuYaRSvsDpSfch6oIr7W8zwYS
9xGfswdn3HR3HEBVecVtnVfOYabP2wZV8AAkHlicAUfIcmPd5qey+rrGc1UMcXEnREwu7F/8EJtm
m9DtyIZaEDKF8HUsToh8B6g/5FXF1zDOOTm++CIOBuwkTePDH51xXtoQWha/PuNPlH5M0DunxYAz
EPvEBUAEc4hW/KDBCWL9x6lm0xP58J/rOXNrtTkF4Jw2uH5pL5IQHyBPspCzUDiQ1JYKhSFS2g42
025kTedQnxymY7N6SEjW8H2rNWINj/HMmo+p38hjeELUZSNSs2SJsv57uY6NqCrMtegOtL3bbMyw
xknJl1gy+VSFTxNOG2DCxh7YPgxnVXeLNf7sMSjCY6QmyGNXERW4A83rSd+ZdQed9cUCEVa5HwTp
E/lHE2eGIMaxbE/1KnV/sYPtAZUyJekWQLz/+qzESavTBixRTnRjEsI1lZwGN7BcRtOYkIENTqWd
iZPZdRFMBBOKuKKKVlpLmlVxu0Do6oTNx6reJpkLqA0AN2IzRHdjYHBT9dGt7tmKf6/pyS8BQkoe
cBqL/V9lD6zUuTmK+hyGPzLi1ec9cOFcYWiK59EiGd3lOPek6YKfl+/Qz4P62js+Jnnft+65Mhlr
sMV7xPAK8QwReOicFV7zUasJzAKj13j2Y8zsaXZIyIoweI+7kavUPnJn2XtSVJT6C84tcKbmxSIx
4FcD+yJE6hQJ3VMn9EG5X3wcit4BFAyJwCXwy4dSNcWd/5RXewBZ5lur3iTWIHw7WGaY70GA3YJQ
dR8Ezufi3DIbJiLGz3uxNKu8nKiwUmFH1hXCpbJlagRCtQWH3bp7dulV1cTm3fglIZyTQUKZ44k/
Dab433xbTugm4Q5WfPY7hSb4dT0gJW+tsawIVKHfYE55DofdvE5+ARPoRDxUyyWsZli8ujVbA8wG
5s+PRS4435e5UYz6PnLqKgYa2eynEnuH3T/V+iBqDLMp9fHa4dgrhw6254xZT4pNMif/h9ruXBiO
eE50zixSE3xiWQ7ZHvb7YzC3ncEtD5FO/VOII01PKX6af0kM95cDWeTI+PmrKzA0FEBqfmrp/QQd
exqOA2jMy+VgZgMMre9nlOgucirTE20X0s4hacl8fbJhQCM6Au6+qH1VFX0h1rOjpOsEdIHxnclK
1ukSUVKFsLGUkGeHSmbASxS+mMFnM3zEBl2OJpr7kyC6TveSDSnwFdUEnyY6Xet04duH6P/k+0Av
SvRTA14sKfSWpRPwRCXRJdq7APLLvq8YLh4gBaV2yH72MhTpiqQwqmsE+kBWpk+SsrqtBb6U4QEa
DnOwVmPs1HsGTwfgmEILnhYCoOTADDPHtMzuH0k2hzM4HAJkaTlZDnVPVz3Ohl+PNqu8aR29GmEc
yKC6VcSXtAXNUnmguW5wy0356nNt6XNyVcKiqLVfOK2LhuIAWw9lf1h+sBZvBS4EU2dMuisF3H5D
fwWIra5XuXY9DVnt4VzlNqboPt6IR2Cr/d4GPCcB/lmDJxe2GRAlHC2xbiocTiPWUwTz5FyvcwD3
x+vwDx3y9/gyy077MRWd4nCSW4qjrVigqtCc+OeI8UvUSHwfv4qQm6sUdUoY74q31fJxveFfuoSg
um1OOaVXcsfk8ks8iKJodbaUHoD9la/L34nj+BMk5/QEaJnOiosmxCsK/QeMxW+d99XJKvpYeo4Q
Hp18inkR5QHoR+u3VJBM/s89b6NQ6Y8htN6PoIL5O18txPg+kAqCNNyfKynKeBIemMPC7SnaqDrm
WDB2+RTQWkhWgQ0rQure5AlZbEvZHCRljMpgFSBEoDIQ1tYA2zWYxr4h4Z0ngJnp7T01A7EE6R9y
B9bZSmgdGHgZ/pt5RyS5txQQW4g6UZiZR9m2tv2vik/5Ve9//KhlicmKJlr6azRusu5i4+ut0HAD
lN2jV6nqD5+z5GKDt8KEzssDSTmuBQg6U+6Cigw0gq75aYM5UTiwP8kjmi4W65ZrZvGN/zEp0TIj
UZ8zima8U8yEqBjiY201liwqf/oYzEEQk4MBTz3TF+mtUyHxXbHumHZvEP4nDhkpG0bT958yT1wl
fhCRZszkfWIi0MBsgbdujN/0rueJQKqDi6QcsMel8KpplKglPP1l91+VJxL/d952tVUr9QNI2UFF
G/yjpQmFTRQj36YwDNyfURQa2Fn/ZJuyzoVXB3l20m5OD44HfOqx9vA8FNk/uqLCccLS48La3nQk
tsNg7p+ElNHzfW5+kRvkEZNRNbg230FJh0fqpXTQyIjisC+N27jodMdFJo3gcjp/mx7Ky9EZ2v9x
qYmWqz4Z5RjBBMR03MGApENc/xgCc6QuFj/xuQOvaijiqPRBhQ5lqLsVqd1DSYmRobbs3Tly5wuP
fMWiUs89VraMQxrvj48O1UvCSDv4rQyHiEWPYWx1UFF3TyZ3SvuXOBJpvvF9hmLkoZhaPBZHZaZj
lSRFnxj/qUCTT6Og9e0CCD1EJHx1iv9HKcTmjz9TG5a6/MfWdQ7IhYTXvPFQVbx7y81zz09PhiWi
9DUTHYTjCtm/2jeV2YY+NhLj/QYu66lj6WFWhO0sLjcNEPhz0mu4mM7HqHxiLBLvY80VDJ4LQeR+
79fJkk8BGsCUVZ9ptzxjFtWIrgoZL2undgxQ4uGkJ0Stvmr88NoZj6TmI0wBWezX3Y0ooDlqvG3K
1smVd8MW8GrSsGc2z2SKiERVcUXIdjzDVgQzj69BYNYKv7PS+ZwAHD7HEGmjwYtrgHP9neVbY4vy
y4djj69d4MmakHvS0HUfCnOVOGtsc2Vs5Ef9jP7emMGue9oiIi1/Hr/KkU9C6DcxTePlEDujlILE
Z8mCWWlFMTlFr8CW3rdYvrmhXHwV6TU4qpjvZ2JzPN3Oh85g0zjbN4dEnQEk6lW4xWXZGk5N97ji
Aa3A9+p01BBNfmklk2zO+Bn5pMZzTo/2RUsTaL/XC4C2OdK5yMxweUHr8qpiQJIZdd/TjrQS2dyd
fcjs0I5ia43viX/M4K+rflenDJBb4U1YBWV2VkzD92jkWzSXrfwDfUmAaR3VodbMsl10TztmKICO
IM2Dv+NS1glqL7Xysol75Klr913Rd8EuP9ja/H1GeK/P0VqWSY6EJp8LXAhlmLupXBrgAV0MSPYl
NoWKlOQJju+Su1I3rNR4pssAWJDmDKCB5UzWD9pboMFdH6GWrRfCc2LG2uqBCAdjMkBy0g5iSigC
rTyauNRt8myyRVQoSZHHD8WpkcvSB35BA4JkxNCe4ndouZ5TVQZdbpJZhB+8Ok2Ux7/HTSVbtyAq
sG46AjLttmt3trmsBDCk1e7TAuYdAGtbN8/FNIoQN76rIBvdkPeeCZSoC919o+jG/Dxkh145uXTZ
xq9nM9MLuyT/KqVXLADLWuwGlT4mLKO32tLXDnkcSkGLIgtHY/5ik5n4pFuemAhkouPcg9cv/tII
c2tFeTtWczJMdIUzmg9x+cTrY3xxZEXXyGpAfwWTCU2ORFuTMshGKbzApUIbIXtSUNa9r31WkCY1
5cLi2PKTv8dRq7UD4vWex6wCEvhPSYUmR8QxQvmqeczvo/4fzcYrmBlcjtqMl9cwRSgWx1dmdKEa
OlIXN97WhAw0Ej09TtBU7+xNfhs8SSZLyXoHrV5FWZNFT+o1DxY9J0rg5bjqOjOpfqArD4mxwDwJ
UoVyxoA8GccXcTFmsn2VHe0VanEn2TJQbjkbDxj1+R1w6WSJTcheU+rslk0IRcI9zaIPCYvuIynO
m4dQ3W7tgFvNR8Iy4WwIJy9VVqX9epNFeS4P5xE9gjg63VioW21QEHuKhnFejRh0o2wmjirOMhNA
IyG4WNS9N73lw+X6NymJvyaFPrj33ZGnDPON1JqxhxDL/3ykChcM35VztErg16GYnLk50Ocee0Kj
YFe7M1+kuOdNUvq+UFi0Nhwnl+IBKN1MC4J9RW6I27as70UoIIuTio08JTZO04F6FP1bCh+W+DjH
FfXyBjseOYyPzrspVD/dq8nZocS5Ab+0Xf9SqJX6KsFdWZBjCmtUqKZAT66bk/DrQ9P2SG62vBql
jlytLzTsfcSaHia9kbKUGfo+u/KyseHCrYgyxF/WEG1Bjbc6/bJo5PSQ60xJEVWAyR+rYvhOLSO4
XVr0JuQ1ScqNvsqdmgVKnH0wkP70qTv8OxDd9yq06PcUHCXdS1k66+AsZPhvDjMmr7eFrHavA85G
96FTSWfn7P2FAJlWnPRwAt2Of/MEwHUGNmrBRGg7lKnBgssRC8imWOEfvsQAVTt4A/sgKDqHD/BI
eaKTgup8D5146KyOhP1iod58aZYjbASoci7AXFCGzh5+eRiTlnA+m3rElg5OmNDpT5pQf4+UHfcO
gPlJJ4goBaXmK5OhxBOiOxsgUFkOS9YI2dYEw2GGkdaq78nYuatq0GbkELdE+qYXNA/OlAy4qJyZ
+WAPU+PzAkc3m2+BSFQf2wkcO5w0r7a6zfRmgglt/GG7OUnlFdFannnO18NIPnczLFORBmRJoIP9
g2TyuDropM2W83Bhk2upjoVq0MxS6HzJ7vRf4TA7IQiG4142ofv39RGDwq1ED2Osab1P55Lc6bHy
U0XDQQ7S3pHmCJ433k4dXvHcxXE3Cwh9D9uSlLYaGNcrGIX7wRsdOQhaY2lcgvhADeEd4hj5WFA1
GaQhhwFcz9o74WdCt5baOmXJap3EKIfI2sJcs3TABC+79slKXJm+8weaL+j5h7duYULafhaxU0pL
k8WpjkXTv+LeyfvQ9tjJj7iBayTBtfLPo6RSN6xifdGLndvmxn+2mMQRnLniQZclsht+cILQdMyz
vEe/iHfw/ojyN8dGrVpdANrDhhv+KEY+/X6FvsMfRK8ZqnLacQcOMaCG6Ici+h29JL9lvgCsvGU3
jWbw5X2teld/6pXIYAZvWQa7pgwzBgZPQoDOP9SD3QLx1rqfVz+Y2zeWIscILePFVuliLHTLc405
7zfXeVgteNtzXdmwguUnppZAilirerYGErl73/XFKPP+dF143HiQVuGD0sPqLMzbA/kyuLrmZwx+
SROj4iBsbat8ei26PT/Ae7DxwVB5v2AXfouSqE67/5jZKt5ZWmPdMWAYpl+5qhSeHJmWJeR+LgAM
1O4uR0zKF3jdB9Pnwp0hDtrUs0jMwmh7tZqGWqHO+QVaCQ0u75CMnwvB2ajUgNf/3YXLLrRa7dVG
5pQrAJgl3myFOnyn7cZjLwbTwtzHt6VVtVktO0BGBjhsWw3zJ/03FtGiRsISt7p/JyeEpq6pnRVf
ilAupOm4HSL1hNAFsuUG9pCANCiOlP5BQ1fR8TF6rm1pZ39j4MsxZtXZp0ahWPgf2M+e80DSeiPu
1Bk/nY2vxmS/MeyWThbMaf0Ro0Eu0aGeHtzvdlfiXfsjngOwYeP19RtLFZX/pXWHq8/Sut5MaKkl
qCYP6satWSy8SutqRKNeWp9KEY+zRHX/cJQt9/fKHE7R2Q5x6wy0c+BFKpEMpy+iSqvJ/Vc+PSUt
eQhwa3JJ1SG9APQptTwlcNAmFqqv3QR7wBsuecAFIUxhnvQp/cU1wpBe4YPtad1vtUkoQPDDuHZw
2zpfqvEvOqcXKYjJLszzrF8Bl3S4xGV+Q9avpfj+tTsxaXn+3w0BzDwGXGs8KgwTnOZpnNPGX7f3
KNnnBsM2vtM0+49uhUpBmuYJ9GfsQKPJTaTU9K3kJWY/grwitF4OqYGZD55Z3BGV2wSKyrOoTxuR
iRKYSciIxEe8bI9PpRXItbZXJKpAjU0eygHrFx65VPIDEKnpzQjydIxyF+pJhhvDvzWf4MDJFuvC
njvcIYwE+c/NSjq42QbMZw5b4paojURjtGkCr/zBAoC7RxIT4vAOL9WQYSFP2N/NujQ9N5tk3z7s
cYXUSxz5UVtoVeSrbgZiGif71QO1DFRfih867KHE3hNgLq4ebn2Fo3Df6m5vZxumhpKJKo1kVJl5
HCw/p3mzHQnmdfdmneDjkJMvUvxiXuY91Qh0lcE/FHOgc1ql353wQeCLB7wBuhL86xD/5r2lYsf3
XugerXOCsSRL/tSNkq9mWpNU3YCwWiCnIqtRTl5C+YZQ09N7WxTFooQeT3SFPIZVCX7s/jZoh/7Y
EcJsSyVWg/qFOSKPwozyWp2vmAffz7cNA33ajNu9lbDzdWYkPkMR2AMQlT7wiwR37mFZ9jZMoras
EkVMwjZgCX2WCf3+rHKIHMCgePAt3a1xAZ/LL9puspZVLbt8QuS5upR6/+ZMBbgfk01Opwn5OMpv
+PeOeVS9ixn6Jrl+mYAQS/K7UEkKN8C36TndoGx+FCA7Y/mowyZLg2r1AqKSRG6FK77vjDQbIvml
Re3aOLTi25VOuaXN/o/Hl3Gb3DsHAARDfXAqrKj3rIRs4Q+lTU5uJLvcESDkoadYbp6QKrs83knD
O20qvJpZtatzP6BAgCtup9aB6QuXm5TN/hkF91DZro7/RKDpGoTGRQlhppcYD1/rWR6NmHqgKi0w
6MBC+FORBVktfpOUPhY+N+dUY4I53v6hKwpyn0p1A5P0NzW96A/4NzAPSyAfYQa9R2P8fzbgeTM2
ulHMiAZ7oYT0UkLIMYu3uoEFpFuY94q2nZMMJoViwwU/fyhDkQMY2GdYRLAmymkvQ1IdVAi4KvxC
wnXtZMSHTv7oS7pVU8YADbcqfeWsfQjBkXvzBs6dDHgyl4qH/guZXXwkx661vKpQM7VH2H5K+gEh
FbcU2B67ORMv+XDT1t+o6b/MQ6d/GllF5Pe399j2zf1ZexU1VNi6e5Tc3MMHVu2/ERL0pvQSZbyk
dRC5tKqNTkTzZCgU4K9X3Rbl6gESTFA9gX9yxfvHF/pcO7C5Zn49lWWkJRFmDe4hXXni9Hn8y3BM
iwR5f7PJl0MOymqp225BJSX9RZK/KtRSeF03Z4ZXjrjGYoCKIQF0vxzQjbRwe22gvB9Zqw0sfBEg
dGMGhEfJw9wApQ77Dg8ysKoWud6FcvEdwSN20EPT075oUwkk3k8eKLAMeUIxcdwbN9S0N5J6sFnF
iZLs9NICouIsd415SXlmeiy07yw2C2MQxqswoLIeJuKmy++UaBd8nD4kxE032F0VLajNROoSDzIf
M6KCqa3YNwtFqD+d542bqaSIx5gwcBv9DsLVY++Iylrqc9CTn5UYMXC5Bpf7wU2ktHiW4Uw30izV
yy2iEJ3yPZaiZLawZCfAVTzJd9fK2FsZa1at/TKaSvYMV+eB8didX1ock7YxEoRneDVsVZtxmKtn
g9NkGfn2765lm+oY8tuQm/7DovAt6T0hDNnSOq2JOJgqw8ambXZnjJpheiQHC02pfSOqMHAsl80L
rGjIQsHrIv8J94WcFd/2e6Src1bQls1WWhBX46RsuVFGKtV2Yx+H25OVsSnrzVP+vsVGldTA2OAv
8P3iDcoojlTQ7B4OyfPfq8qlhKGn55azaW+GwI/Jg30GnD8w9EB0zF4m7zRzXXFAIKEm9A8LiGhM
9TZyqO+grGtnXTXepPchyt3nkti9AtjKIhc6ZIEjZVOy8cjAHzMkzjEk4Gn7C7sJNXCqgqkDVCLm
1xlzvkw+WiwDk+/KzL8tqbb2K5m+WbYi4xOYK7P8qdkhzZwxbkuRYTYBWEK7UIzls9D7Yx3Vogbf
YVDpDpVGXJg4/drf37ZwRVfEzBvUDEs4qOnJ6pQE3FesGAIAYLddPgUeN9eGlfE9SYfZwaQkjsYO
YdIp2ytM9RbX9HU3bMPwHhQ9sYMvWRjmtVGSeyacHkuhAGe5touF7mFo+vzHWZ41TtBtI9+8BrKr
Ba4629yrAMt4uJRYkoPEz4fUNysfpoE/TRKajQ6hCdBFNzAGT/FgJ+GoHcXw0ZgXqUDkQmEX0Uiq
0W5helwrv5YF2mLQWGLOAdvQBCelZIjYU5Iv931i3EKfROs3IddOtuJH+IPMa0zFWH79/8ihFniy
VbwCoNKj8pB/BlkLDVLG+Fcm/MSzlsiyyLfE68ve9zc6ltqLsWi0xY7lLI3ad30NF3Ox8zmkgM0I
XLcv7ihFfjIJER0+54HwhtzUFyQdXLHx/1/AEpe1Ar1Tzt8wyhCFJH110us7v1o4i8k7uuKkjOob
nt7GqWKXXOxAVmBGYlmLjWHrXa9F/PXWelCR1MnBF2BZjNHbs/A9vNeQNLYWBYR2KxWiI7v8JvmV
X+rqoaRE1uQpdojF5aee3tEYb1FnJqycIK+HNkRkteT1YNEpUeGEhiUde+s4KS6YM3Y2ZLGPJPQO
udER7HWY4zmt7eLqdRFBJCvHbGDnBI3YqLB/saprhCmE8r3hWdJgZESTb9ny2CAlCWIlcyXuZ8cB
4soTedCHMkdqI5KejdpQAsHdS5/zYgeri74kDp/rSgjRU+9yXL72wfQRrkuDF8i/shfgXgODW1A0
h6rSl/921QhUh6oqekRMjl9d/eb2dCPnuYLSR8WM5D3qBj7qoLBgOD5bNDJA8vRt3V/bzI1Uoi4f
Rrv4xcoczaAqLIQOpLDGfvbBxFOs/JhruImOJkmPcRGpsJosZ/QnjunuRDWA1Pd25OSCv7FHwOKM
fL2JWd9wdy9l0J6BrRUe+y8+qBZcPZKkA9S/UH81D7zl/5I19fELpKGXkvsIJ/SPCpT3OYbopbcd
2RNUbkgXJlB8UA8EyrQfBgbDAHPN4yx3KbS7cL9m28e/CAJ8t234V6KHoqLMNotbw44gPK8qtwMc
Sn3FK783Yp5J+E2DmYbTibmrTBMijGKO+fDnxh4xpzpjBxwgiExl9BOtk/PfNmDx++9zg4zyr87M
v+2uJ3ZA/1g+QsmziH5IpOP9A5Ooryze+JlFuKltsBMS5t8+1Cw6sf3SSKxCW1JoJ5go8iyHMKPx
MI5UWF2/159mKDk3GlHt7vXd3sW6EhC+7CfAWDHBy/JWUIRnTIRkxKaq7WWmzwJcp4AnS62UAT93
n82EvZY1HjXUceZVPJdpSNrJaAZppsAxLOiHUDMMORGZypMbzEUtI57fclhcJXhU+JHKWXy9c+vW
hgOpJRP6CMaLDnSUSOJnK3mysgl16PIaeg6BaZbeu9UfhpsU6Rmb1GnPxQzZtpt3WdNvf36Cpi2f
mLIG84fgv5pm4Eo1LOhK8OJ4iSVsbAEZQBbOQeY+g13T1UfygH9mJ4JDS1/ijQYRfXJmCotju6NQ
CfzcSqXK5iPGk1s7KyturbjGBevordmu7YBG9CT3Ne6w8mAINl5F93DYfmDsjwhQCvGLs+q5Kozf
eBuNVCDCLn/pXXFcqV87P5qubKlSFC2GPKF1PhvZcWQrmF7+z/kaXmeben1JWAU48WxLbnK/5jWJ
T8FqDt4iW2v2t/ll6pdfpIUS079YNFPxLdDQrOk++wTw9i9dg/co9gOsffFALchz9h23+3IAaeqZ
0VRk88syeW5kYCOePeQN92ipO0gdLfK7mQenoGeS86yPFtlFv+4g3a0UZTPgifUXaQUWyd41gocy
vhwqEFDOUHLbnNaqgLPUPFq1UGOvIgq1gBxQfOAK/XywK8NShgir3KONEvjmKU2vxmyo5JI9wvGP
oUheCGNC2Sq0wMD5SgPYDeXt3ldXDeE6pT/N4gmRVd0l6jNIU5DMf4+jipOdkzJ/usdElUw/R1G+
YdfCYgeixBsBfx0PIBSwMGZm/nM7x0iaeKxTGbqxA9FWlafL6rml5C3O6DixVW9Yf8PH20bX4wRK
C+dXpPsLFGuyaiHboABLQJl2YpcFBvOfw0wAMNfqESRw5BGLehIY6pi2F3K3mnZ1k5dJP4FASjOT
+EAc2mpzxWXQcsJeERU3sdskqrydYVOX8rOowXS1u8ShNjZMVC5OOZt1FFm+njDXCsYkXs0foEV/
1bxnyxqzww5F2WUwnkkXpLQ0jDZaqUDw/jVaKNGbge59cyj6BNd1qllVZ76q0GfSHHp9nTGjvTYf
6NHtoYFJB1p02IOkNPwGxBu6iGZNH/SMtqejTBnwESLQqvRij6Rg4hRufAob0/MzdAwmdbgDh4DA
9Q9GPZVH+Y3GiJxuRQIfkuwTeI1QTCIQNKurBMrFJhF1udRcw6rpxQAQwIx+3AuC7QDAkQ0VkH5X
MAXWTF35QqREggYfCpcbvJ84z+4Z8zl47ZG80xWubyjxNVb6PqAF7HYXOfx4BroZz35+rjR3JuUJ
TePM6VW16v0qIgPBD5KvwTj3ecAA4ISCH5cBH2awUYR1FTpAAsBhjHw1sB2FuUH8/bcaLc2w04GV
gHiYXb9T8aJ2zpd7C5fkCUJvrBCDpXIxVaKoisCszWhrJxNu+G4lub20I8ZbarjZgcZ4WVc/Evm6
+ZoyvEuVdfRhQHqrz6D1nUGdBIZCu6KAFmNKoj/OgqQFpBvhxlFYvgQBzQtB2+urrjmd5hgBeiO7
Asp/uRlHXsxLuBSWs0mxmnUXIHgCMJYK0xoVcEeJ2tTOEaEFXFoBa4m1gE2M4L4DTqegNB6b+I99
UaWYazSFLhbYysIhFEjL97OqqbCDBrGVyGE+jrjHZPG6s5v2qk+FeagfwyQjoFF9GAcBuZ5L/SS1
9vpppoTRulmXSqzrE9f0wEJec5ohLVObep9ZX3RXUqDUChkcCIEI5V8ixPlrjPDfkEAP3BGpRBnM
otNu2QiJCSg8gOmp0Wsbaba4AQ+XGiKna68gnOqb+MfE/X126K6A4HV6xe81eFgGdz7wm8DiYgSY
FPWgpJU08zV/rVLUsbMzFZzQp38DfFEGmUYLjM7L+OG4cdkRExoi8aMr0TiSK0Cv2ccbwJHylKFZ
o3NhrGR4rYg/uyaCNzblaRJEtFQF9jShFjQSpOXhZkqwntbQeWMPoQRkZV/R4/eubxKMR6qM7Hs1
NvHnLnbi73NxBipxeAa8TmgS+/vnuAr6w+eN2wfDXFeqZm+HHU2exYMaxOD6jgSVzEJW8MnV35gq
r9RDiroyXmI/t1sn6zRmasdSn+YYIPB4QUe/evVZCjjTahownWuAPpyRkxgNI+XCXbwrjV01HY8c
Bt2cvTdJzztwQeHrfWFsYSKNK3LycYLm06KBvNKkT5WzQqud2otRRarTkMGMEcGD3XxOHaePxXHt
m9K4f6YPjz/3y9CsXvbJ/n9RDbyouz8FnMw8XCgUHI6bMBjtdJAcoSbhUVcpXMXE60Xz4bpJLDPF
9LUbRmz1KLct0KNI1HEq+BvCVTKd4eNberMyI0KkVhCBo9nyVABgy210GJGDDAiCd/3AeJX0mMaQ
kYHFwCck1PROoFxvBYi0DucGyl58PxU+22n/a/FHcY55CuIDm6rU5gLtmopG+c//pvwT0gLfbfbr
L/gY3P8ber3EvtcX2p7Q5nEOTWMVWxBiDJ2PycGIzxINFGmdpiYjG7MHdWqYlisvABY3JI3LU0Yc
2rBLQapT3iPmWH4B9Q2WV1E9BGqTmZ5uhOcE+a9eSID61gpFXYKrY5Cdm1Z8wIDh2DJCNnkFvXZz
xXQwomsu0ILW/SeMrnHhXXTuniTs4mMmXt+Bbm9MOoZIh9KRSX1/WiSB6X2fe82Bqrf9olACN/QO
ySIgO0ajLirDaSFiRvW65cgZtSySe3ScPeA6l7gTi5Qey3RKMI5nm0cZv0pqqHw1uDoM1VuWmkfD
b7Rb09kPUGNLR68RWC+vyulNKYsNNnTsG6WRUTSuPHieMFLCvq0lODeDqaXJH1ICEdc4LPbbv+u3
YJQ2sJg4OfFigtJeShmKaObxeE6uTJvIEF0xWGjMw7ACdWAwIHak6i7uupJ9zZrdD0RUO2Il2Mhj
kd18WlSk+tDu4zX2JPwuC0dmCvUAt1VZ9jQROs6GermP1hsMKeYDDURpsou/enM7mU7rxPJBPWpP
TbnNejxtox4VdhywQdmgpl3iSWtozl3fDi3oFNFAbNGc6X5hKUqy8mMc6BLGdGscdhB7rfnxHHsr
YGuK8RkVxXirhAO7zhLlEevvcgQcEaJ+6Iw3Zok9HHy4bqUbczXRWWN/8+6J/svQFEvnI2jOY7gD
i+gN08KNoEsp0VySE1CY1fKP/3RfPZJTKoBpGLIpYjP5tzIIIxe9EETzzTSaI8jmrF3jN1sdTPT0
BQt9KjBC5JXeSCnJSbPvVAKnMCiJHlqmtYuoMlODo1RTb9Wvskvk6Oe3HXCjX6ItmQ2Uap68vEZD
dPHuNSk+0ZJQCuyDyZM2Hwe1lK/ipbFu3icTY9ydiNG88kvFLrRPGQ2UzJjF+WI/YEXG+O9hq9yy
Wc6xKotQCN46k+AZzBTR5Z1ouADRBKsxVgC//VKQSmwTcEey415FLFk5/7YL03lsnZvteq8wvTo6
UbQt+HnPyTzLayy66lK/ZH0mG2aJ5pec/O4M83p3kBEHMaPw2RLDjpgZHbMkZEaPAqnCBVlYwbqX
n14KIgsLBCzfIzoIfR2LoMuVQ3QZlcE4PLIj+2ySiuHYBsMH9xpDrXGVu/yyJ28WVaKn/xY+QeKD
0N7wJZKggQ0SdcccA9+Cp1TU3EVoN0UvhNr6Lu7If5LeiWCUpRzxD9HFnlDVbMBZPGbG6lqZU0Sw
PWY9HyRQYpyX3pQxE08VWVi5mmVZxovll8DmZYUhL0vM6waGUXKrGbGfK+h3UibSb3wwWSoCHjkh
Nyn53fzKMtEfcx3iyeFl+T+kOvZnFce/TGA3+s0H30JFp6pAGWGeh6/yh6Q/VoOYS/BoGpfEVyTk
I/VGKTlBod7ZIN0uA8i/7WoPZWTOKOCxLHgtMh3nDVq5ST8M3QiheNl9NhP8Wra5n/eJDRck9+L0
GZzpIvYZh7+NGWpQgxa3zyVrNRwEX/CFKFAckcHvz6MHCmQe5+5poYWGFdtnu3Ci2ATJrxA20u5H
XYrRmzFdDVJ50W74e0oBy31mtcaPKybXw8aCFzrU1P4qHvJOhe18Fp21AuKFUyhCxMWpoirbep7n
rTUVEOvqc7VYy0L7qLWGCNU2EHfDKgTh0O+osFk/b0NgaOjzA+YaSMf1Z6wk5WXjgFuh4hv1e9kb
kd/moe5Q/eamtvaB7wHVE9aos/b45Kr+gX+3PeI/HOaFEnpRwX9Ms555i/MPGWHfZ5UoU/VE1XpE
St2tnRx9+RjqKnYZVlb48n5jwIji6WfKZn010wMOoyuCV2kREoLBE/VHfRiKHnQJ9DFSUx5U/9Sx
ehzpnDCzrTdSqqa9+PsPLoczpdyZwboeZHflK0Dkmwm+iV9AnLa3AphhgL4prfp8c6o9oOoXlqTt
fxye7c6yHHjRRYLtzdZCWV0JWjGlxaa+tgQPOrXIWzRjMdXwADcUGcu9yhwoMQMApRve/7u3FpF4
YY9dSPKUL1iAQGVgpL5sBWtmtyhUZKR/Xk4zRHY6EiYDhz5eYdCGt+zghujfXVtS9iZzXglwa9fH
VAR2qST+yHv/Rzw3+YtIiCYuemki78xudMfs1BKrCrHAotj3jweLmOG3hm57EqPQvw+CGniv1VLe
WE1v4XanlyT3n+N+xTY2pqi0lWlmyIJ4iflOLRxc++VxANa4LD96AkV+v6luxEPRXWhMhKJpKvmF
m6UcUpmBHb3KgKmVMvwIpPBkOBIYgRcdn9iUUOm5CwRxuNpxabjW66A4vMS0K1iEvaz6d0vpexpj
JwJ8+MbOFRLAxEWcYyqqZVX1pb2f/N3d2B3TNNT+1SNpBfXS0Di3m0tCcvfiZdA1pSywZyqRj2CT
PAe0lLuQdIKqlNAC0Rs37Speu4Cf3gRgBCIBrtqtr9Px+Jtvk4M40F5+pANSCzUwPYgo12klB5Tg
Aq18oeCbLhkCPXmQdh2vsM5uvJSednYs4RQX3I9heeNUwYFejf/BmT50Z1GdWrp/Gm8y8Nb7AuO8
ZKklyRp1rjiRcuL++ioraK+SsXm1qnhhwGqJrfXgh842t8hLtXoe+n0TbnSYeSy4ofp3uV47p3fI
LtVaP0LzaCiaMMN2jZqmL1KYG72eYxBEeluja4sbSET0OA9h/g4drY08K1KfCbJ29d/AD2vB9xvp
3r6d0kk1qp6ychCV1hBnACmPdkXiXLyl+abA4snOXWCPIzDW7ec+b8Pn1NV5Xu2LRfd9vJ2bAEcM
2iz7nHlTMYeH/k3FgyufQnnjZov8VGJ45DmG5yOJWog8ULQqWzXOr+dBru0u2tgUbD+0g7LRJhqJ
oJhOWi2atVDnc/MfojJR7yZrg4a1SHqEsV53r0yVZr9LIZ8WNWPyHCXx83khREi05dEP59ncmmNZ
yv65P86S0A4q9klyogaC27AxDMbRDTe6buYutxcuEjqLW+yn0Qb57XfTY1Ekd1BR6ihNO4I8ZPc0
nhfS7gImUJObGouxRfenTm1AIx3arU90JXf5QCbE6FFvmCKntw6WhRYoKarDGgALddFniaAweHzh
zZ4d4UhwYbajAg1cm9wX4YVh+4aiLeK9ML+iezIDMr+qHx304Ezp6f31yldH9sOx4ArfJN0Arbmk
R26kA/PsUHNnX+9ZJJ4OiZ/uXY3nWH9v/a7wUFEIP/FPEIPViLJIzmZliB753tp9ZIRlE1xBgbIJ
IhhbKqSZJclt6iLjYJL8W1vMu1ck7rf5ILwrs05it0vIEdPO73cjH0cRgXdUnqJ/oRYTHtC8ZlgA
GCPCdtxmOcOUH0ibRDPP7uiGbZ9I4XVjGSlhi+FVMyPgZow4tqXdKJ1ecs3KVpc59WdURYcEJdi9
PDYPIVaWEsbsWdI7AFTD2vPKZPIsEDPsoKUvPeBNyBzzKMCbehFV5PqZYQUe9VFQBP2Me2w4eW6w
o2bi2jPpefwJV59tfmpo5lYfHIN6u5PZh9m5Wu5xwbeB/quIv1wIXShnEKIRuAfNU7qhiH8A1DsS
7GElhOUgnK0QeEP/X9zEX+2Ym3SfT4+dsBkHYWMadJrp/bGxdAa6VDDYUJmynVbeoA7tmxN4d3zG
jdeiGw5KPLMoh3Q62AVsAdYIpcOUxIbDWqWQmmk8ExY5kUhE7wpj/RLm39LFdBEiIGr1dqjyhE3m
a+PHit/RfWPtywk4rXUmjnknx5ThP1r2MKD8Y2AZWShgseJGRvxrwJZiB974/P0B5K2Tqt8+Z4ak
weplDXxbtYixOKkm+Kc6gZiY4075L8IHyCyWzY5obcYwtm2YFPp7y8SiEZjONfgu+vcS4CNwEDEp
3JhY2sizQ57jEl1XpsIG7Xvpwoz6r9pNUWR8ndb/rMJNJm/bAbhgMy7JJVlyUrC91hjRr6Dqy+1j
4uVDqcTkkBBoVdvIMUcCUCi3bi5qyB8GxCfoTIl8LAYa7MewdZWgkpy83g8gNZwi2BUvC0z4D/0x
QrpNasvWLaIgoac04qKt53KJ3zoAR2c6WLwx1bDCREupHmcM+8wx4ogTt6UZnFc6BuiMNEYPI1Md
pjxs4/PBUcNm8sZEtPuPzPc3hG9qV+X3mBjNqpqcH+n8F8Sb7yrnLojtN724T9l5bsbyXEmxyphW
O8e6MAhagzymBWuOy+eUvJc7dGzbTk4wYkjxlQBJ3mw82Lxgr2wIb4V63Q9yQieurWCBHD/vuoMw
63YNjRMaSGChA6nqTDLW7O0yvvw7BupnIdI53W82yAflahwRQoNd/RiVkvPub/7rpzHA6wSfuPu9
ggTkD34QrKaO+XjxksKnrNmBMXhA1mX4Mk3n7GEW2/CuhnbwJRVsRchE/TGKqlSLX7jM60ZZFfea
0jRsQ+Wzwxd4Bfl4tvx6mPXm3LpM4HJgJQpSOUxKhwHkj2j562u2NKV+bC9A/iwuQblQKAPitW3E
+smlk/Wyd9o/nO7je1Oep4HqQukRWIsOPvpsoetCnbtALm2rpwJBlKSs47krYN+QOe7yJf+nE61v
xaVvuFoerZyCBSecldMFGKmUlxwN3eOK+XkwVN6UnE0ybDH2sCDFb5woaEo523u3w3RcdwqKZjS2
z/XKK4r4UPJhcFTOd7NdPveCZ2HnzsDkA57qTj9NfMgshBy2KSSH7RmYKyeM/i9wIYZOlMCgHjnZ
+V764SJbN/6aUVrl6Mf9wy+ePYTHTP2YTEnhMRS6tRRoENoRY9CPLITykXhc+Una/abOvmzvHJsJ
iySVWL0qByIguaB9rdAgIn/Sq1ra1NvrhZrnSv7QfIEXHY/NadKE8JsIzATpzu8VTqvMXjw3QnAF
H1r3Y97hD4+p17/SzAThWj5AXb3pzkcUz5JFG4KTL7cn8TaqN1MPbP6ISb7g6fOq3bn+JRfiMUQp
/XGcSd1Uk+JHbDEPzLwSOtC6wZ/C1GuflH55OiG7CtH4+Gvj8bR37/KscU/3+USHJj/mRgm8GbJt
wjKR0swj4aboUJBbF4mo6LYwQcXj8NwbmE8+A1mjP+NBaPZwZR2G4VOxEtKnGPhpFqxXv+0D0Gzj
kIPqSoO4yu9dzyjbktfRJsTrwPVgtwduq3RiwZ9ySxA1u6/D3D3C9b5wS7lxHmNtt8iv6GeK5IPV
Zm20R3Eb0N3wcc2LnScJdT8NpgZvoGes1qPngc0131ak7mJBgksM+JsQleNoyRXxXZOCrrRNvKYC
q45d+7gq1tDjguG74dCKzZDVh6/8Tk/gIf9rJ6SnXA+sv9hCzezw+9x16OWjCZgArgjYsgznW7OH
X5eSZcdREOuj6HcgpzfZjrD4+fWUaixbs+V9ddUllG8sWNdTYekm/c8E79mFsUSAbY+QQnNljLEQ
KbzaDLyBHO4ScxHnGXAE/NubOThsy2afLFgWghKRu9oY1jvdie/A6Lx9Li54l/yIfDXTK3ckX67q
EaDM1ZIwqOEq4kpSS7Cchtt3qVUvForozyxZyMNJOa1ew2N8s8nSXeMvko8mBr/rtDB9yt1JK2b6
tkqyP6DDAyPqrN/A6Hfvvtt2Z4v3kdqkpE+H5bBJmaWV8Y8BlQgAvS/2Ak1qSfwnM0aU9mkWPW2c
hGlz7bwvVGAxFSFEkuOQayf36xPcD4sVs2YPxdOAzEqJXIIioXTNY+VBf5p4ZNYw37enEQM40sR9
pKWmOC2Kq8f5eGrXrs4+/2hmGX2T6EivIpaBwT1dYrsKcrhTp4EJnnf24LdNVuqL2HYQ0wi5fv2Y
5XmZIToxd96aChaAv8CYShZSq2W6kmeSpgMdItO1/IeizS2Oarww0JxTvBOEvnt8kKGfKw9Yb836
xD04CQkXHIWS0wEgI9GoadurvDTk9C9++BWs67tw6hwFO+E3N+VPycDtsF+wg1FpfqqpYpHb3esM
PN4dpFyzA2VwXjxDVbu1eyzFLdzDxspFemwaHFV+kbIFAx+u7th5foBu8PWkOE2tBP4TV8DnjkH+
9OcFNLwp7eA8hr5LprAoiQjw3A6clo0FMvmkFig714zd7vDwZSYVr1THOijFPYb+016oyGkVm7/m
pg3HTY+A7+7csyc2bvbAEMBFBoOptgcFpf5EEMWvd1mrXQZlXHuyT3QTXY0qcUAwdPilTK9qBFJX
qABNXbcMhUnzDw6+WgfB1cRZjmkuw7PV5uR01JXubR0VRIqrf8ZYmqvOU89drRgMKhT2zGDPJtjm
oU+CyZFeykPC/8pmhTLfDyNQl2YrhnNu8dPPERJuT6wxI2/VGia5DNNQrQgj0k3XYRAoXf38dcvN
pPimnkV7I3T2NmMaKFJdqgjA0/KJERUPY+5IQxAFoZO7tpIt+J9vjyWlkgP0XbJZRPtEOscRHTNb
d2PjgSbspchCkrt+QPrKFMXkscg+DUPhgO/RFaQh7bOlmxQTlO3oVOXPOElHemjA/3Ol36dFjVOm
cJBqslTMwkDpaaF/wgnot9P+LTasPjW1bvsrJLjtT5mqOFGqBbvmh5EvYMwgT7qbzyAMQ4Ny2qPi
g3kbL3Uz1tR7LVE2gR/cR9KFRrfuo/2UlZ9Zw+i3Vnv3gJ2azH4sjRQvS8gDiuMk1pj6b+i9IcCY
yv5jMwSdwvRDoAb0RjzLVG1Q0DacjRmpKxHZXJpuruEkyrQz66NPKWdoSTwrkONB9k5m+z//eQtz
AJuRUWTF+EqD94vxIVf/0O5JNG15iQxVTAuT4d8w4Nvf5Bva3Vn9DehjCv3e8uQx7PrsugX4p/cN
QsSQoml0FX1vIQxjbqpgjcZKVvKb9lNgnltE1rQzj8E/qSQZmydN8hhhavotjOf4nAh3tW4cqlc4
2PWyJUPnFBKXPSOdd9gd0GAkWTtIJNnM20JziRuTYVtH67hLHiYPEhoeo7VBiBX+YnX2FycXoRu9
EFtIla0DJ3JUXFBpEl3qEEG3SqirUaGdvY3WvEdcUXHpEcsIxxsEVd96Jk789flcstBxR+LtEYHG
Yqs1AcPP1l+Uq0kNRnRJMCxIL1wPhXKiQqtD5rygVKEm2lhogvg/fEOJgJc3MTGXfegmPpcwCVp2
3MwXqVpVeF2mbnSlrGi+iivgGmVtlPoqAZQ+jA9Yiypa4iVE8TAXvpa3UA0B7CwJxzY64h8xU6PM
++VCkBLjvtAIWGsLE2qBs9SkdVkb0TpCeCN/udctmZ9RlSphgfn1avEQ6a3GNFngkUeNbWIvLdNq
C97/SYIiZijFgxaC2vavGb/4XmLKb657YiBw8sRrGRfAgPhTh0ggwL1MDPXLQkuzpySCYa859VOh
u0DbtAKcVlS7xtyfLzmclBp09SrCKQ1Unopggv6WR+nXbMuho8bjC63oDS/qQiA/EVukdtnwCFOl
XZn8p6ubYc9gSN2I3/uNQlDgmsC5zq1z5nDlW/g7cYYjm2c0NrEo5oPJfuT6vd1e+XMDiStMB/j8
j93vNxeK1bJ/mO3uwrOHwFjDbJ0ieHiNsuTh3ViVfhk8O2C2zuk8lKZyKVTNhgW63YGOyBqhpGIv
8+xvLdyA4KprKi75oJd1h9VP0gSkrVCLbzJS9ZFWUm12K5/kyzLQM/zfsrq9dKqz6+6ZAuWAACDX
62xxgO7kaBwE9lA5y4xHKgQFTvWhVv+5zPYekRQrcDJx+M70nSmd1QAV9CfxaJO76WJbor9g4BA7
7138Roez2bKG5DXySqJ/w4vHtnr3RrjIU4+ujM63gfc2T28STzFJbJwYKHhrTrxLEgP47rZ+DKd8
+K3souIwVe4I2NnmfXRxiHJb1AMackkhQMb/m+lFlEE4phUZlyk/e9DLjhV8SeFfHR6Z19EJdHPN
3OabknWSXYc03jvpP7wWqccDWMy7i1EELUo4Awd4eD1B5b4Zi773TbqmnyV899Rv0N6gFuO6kWzz
nHXpHE+xjMFdMme5eM5CdXLKmH0tSfAm2bo1I3BcuFCZ0ki4L/tlocPDWrvdzbI/EtOnIKrnsw+d
QBIFhRwR7b2GL9204R1jJP4qNfwuLaIGsRr250a3q2tZWW8ag6NygI8qIYlY8bqHJGVUDIsZWA1M
y+LR+twnQhPYezf/oOwfaK7ErIwsD0Fr6uYh05B79J8JBKKz5nqB1RjzaxAyOgfQwrYfQkYidc29
+GcztEn25wwLKEoiTjqi6hojQbxVFq43NKc3ipyiggUPDFrDfr2UwVu4Lyd4bSp23yi2zsRBP07v
Vz6YV9CJ+B5K7WCCD2JKAR0th1kHytnkH1OeZHMQj3bDZuayUvIrIhlGMm78OznpNKD3AxmufKzQ
lrWBe+I4kgKcGA6MK7lTUp1+SY+tFQTnX0b8CjASb41zMW0yKO6SlWAk5EE0LDg68pIRZasXKZNP
iLcFJDM0H1/GTkcucOwc/x3kfKLSbFHCSb/iPp22VQI3V+hiXiL0p7KVlrIrWXp7SxDLDsiYiF27
NiSzeVyl+B0JBXkgz7zSs3zBICufzMYrgID4bdf8ub9EUqUHI5SLJ2rvuNmIVVbNrVpmDOTrfM72
bFL0RA44JKmXJD3iHttTUfoNmG23erhCd4nVqEbvIg0zzt1LDYTByaXPJqTrm/ltG1TYQWYrHegE
T2Mg73JAO9LsIdFFEF1apf5ZxAEIqcyeexJIMvtMmHKw9bAVcb3eXol/aXcPOM/fiQnASegfAEvZ
xm1Fnok4kvAkLkTA0PeIl06zU4In1JwEA83dJH1MlyZG1H+8XyQmQ2WPlT+zXZaDCcOQC8Ye6Km5
L+KQILEmni2RUCWGkhCF1k4XIeiAPRRVlBkvO81f3HoUhF4qGlei45yHYNG8sMtEX6O44v627PXa
PSJ+yxe1tbZD6+CqhRVhZJnahqYXBO88CeEiIJlx175866xuH2WJc8c9lUavbIxk+GXEliDLlw2o
hc46N00s78Fyvm/7K0w7+v0QzsSAQ5bkVeBQ8sA24Id8XiiLnmNXudthHUEsywDkCcEsZIAyf1od
ntwJWnXOca2CVUenOmMPpE46K4G0ADXl4lbkRBqdTpyfJ4oToVXWOE49/bx8GqFvOyUuiSuaezbK
ol+vZ/5DPdKvVFBszKCpavJsSXnh/OO1BkA8UtN2lDJQJtXuZCvWMX8HAcAl/VRu3B6erDQ+l6FX
rh6cTdet6CVMuCcon8Wjo/68MBAA+WcG1k9F/PBN/uHJx5v52I6sJdY7HvauviSt246HA5hYNlsf
N0oU9MKp8POOW2nqDoTeFaxjSu4b6IBFy26KAIq5pWZO28sLmeKSOw9IOQcSMGg+dfIbHk9P7R/X
XMByl1y9+0BNbRL/1Oc1dNDvGMA+1yVn9g2neL647o3nhLC2lQ6O1g1pyRQALqALdFeirwMg4KdV
rvyDiS5ppT402xgR7PANqnL75SzaFmerSK6XIMmdyySypl1u2WDIP82oGW6/O5Wd36zzDTCzdDA0
JB5BRFvLLYQ6PzYH1Fx5aXDnMnNbytoblbeYNrOfQZR+k6/vZQbI5hIVTp7idWNxFNqjsaliGZ+9
54YSjVo4j30apTcHrHAXAa6oty5A8OYyL2aVZ83hhb/maGN9egslOPQQjZ4Seym4Cts0GLOv4Zvv
LCDPNYn7HBMXObnv/gIGuHX0CsSxN3cY+bLEPZ+QeO6LFFCASolRIJgYChdkFdgltrt680EIUJvU
xW5Lq/ZTuZUOquXu8JUi4nLMcT2RLdMxxMIE9GGFmE3SNyObmdFihhldui3C0IDIGAcvSOwzZDji
+7VCHdZXUAEIdizynkuZmw6T/Xx1xCiTRd95+y0vvSbsel823c7VQxQOgwgXv/x2ocVUSmjdVhrO
WwvDRQAnq6N5BzrZ54DVSsP0fosrXBeen4Ro6MQEeM78HTsIMV7pEAHlK8JovzaNiDfL7hb0MojH
n1czCzI+pXymRavIocuMLH/1T4WiPR6o5gKxiMOjS+7e17/p1PFydJoS2DMFM3ApyRqb7VkIBkFI
SEPgGghVS7XDe277o+9/9s3AfBe2aVRtWHC6ikqzBNkeWNqrXjR4R9/Q3Fj4FRC9v3zLoAC5dSC2
z1XHBWbAPmC397W8c862qUymJYKon9k99bv8qV8XCM2YTbZ+lhJo4xp6AX8CP3SJTHENUUnMKy36
K+LIJTQB5nySyxzBpRR+7cJ86Vl0Mqy4Z2Ihff6lxeVt5i1OE1GN9O5Lfj6qyZFFMLeXIXgN/J4k
e/Ae/gUK5eTM/eogRROUmn/33CccPtjZANzR6EcQTpy0rLF66OOOg7qgbQ70QBuXU9Z2cYYn1CzH
R9QMDPf1crD9ci3aLy8Pb5bB4a8r4cuItHTr3HHegAiEP5hD+eSL7H4g9rrd8yuzTllmZYA+zu/3
u2kN8GZFvn83HgLQIrrs+mXwANFXsbK5t7uc3UEllBpb1kRd2/tHMlDImDbh/rE8XWNb4Fm/Vd2r
J8tNftLKwn8mGVBDoFp44RSqQbD41JEhpkYfRnVdE0111k0zHMjHXphV1j7CEQtBdbyYjFx1k+kM
9N3FCFj2PrfnOLeBR8ra5Xv+h6RC9hLvVMEQXC/k1cq/RTg6WsxavBhG/pmcnRXHhgKLrOS7Mlp3
vyAtOzLQ4KLzBlH7e/hMz1EWKvw5gOYhkLJ0prvYwNq6ofVJ/nWFqZTMSun3eXRnaOVCoNkar+Hv
V6xw+tZKTd9PW54skbwUR1foG6YSucmjasFlIEyd2k6FxIAY8GWnfo80u+a9GHXyB9ycRF1EsFjm
IMO0p80i1IG/EMKHMVQNHIlCVFS3NU1IdOXdJD8UoZd3u452pfL974y7vmVzKCL9xVIpTrhzQPMD
1R7virI9rRpQ/RuKeXJjaPNKMXRFMb8bloiHzMVQMB34oP82IVZ/1UnemNtoRSwhhJSm9CngP7kN
8iLsxfKA4MaIy/ByAGWwA0FghPM+N7vgDy1XHA4f0tFtqglvqT21bEfUHB3ojdse6XxTC1cOMkni
IVmsCyhkesPoT6/s4ZdXKgBIWE4w0x/PdHqigEC7JCYIqUWJ1Y79xFaorWsR8qr6a5W+F6CV/D4t
i4C/erdNzw9XLoSAR7Qe435BzRGrVqQfV0FdvSybdQ9ua1oXXA0DdnT5Hhs9J68vE0swul32lmIE
umvVj0CiMvW5QNLCnlLBv8HpAD1WlsduTuqFvmhSl/P2GdjsmbmMz1lvA55qlKFm5JPkZE09RSfS
RNfH9CTPfoxT5Yp1l8g49lEsKXfybm06XjAUHM6rrch1D5ZeupgKRAmtzL8YV4yvu53RlWqR5Pe6
VVoX8LeMCjJfiqnv6+RsL8axtO9b9iRBiK17CbLCeiVryTIMF9aAVgMbxJLFk1gKCMpRdPDq2G+z
SRURtdBLZPZzYbwx5CwOtY2GrwRg/z9tMIx/md0YysAP1+Kl4YdGk39mOGoWFqBC3gw32XoHvSRJ
TXywHfbnC9vH6Bx4+xH21qEbuPXutBNufbRyl3ePdflCZKQu/KagmNgd3nPVHWms0+qyHcFS/nFQ
j/PBZBGKfQ3smDpZi6RP4/ZU3MGi1oeRVYadzZ4MFVZriekDz5jCOuZhhTsH3bwk4wyPzrHhNSh7
dZF5mNhtr5PkJS9z70Qj29YxhEOUHJX51Mhvk4+cDV5nyqRaZBunysPhd3TxQH90cdcUFgTxKRBR
fw0U+JzNfb6a4VlsTuJDXYam1PMxG/2K6hNkFtr6YftLH3L4xH5Kt791qX4Bj8U1cY1XqRCYSKM1
BgMo5L+n8DDocbQNFdopTAp1VlvTx99Xcsouo1pPS2KsJydEWzlDReHW2raBfJbQJ/gKzM+/xpmo
qZtPeEcfGPcyjffcbK3rPJaMv6ILhB7HL+tTv50GAxSAbQ8fOCFn+Kg95sSPAF85dNZQ5q5j/IEY
04LtcddGnltO2HU9DpmLek96znFL3dVmE11Lsz0Rmwk178bi+yrrvO0IekbBIoqtA+5Q5oQHVI0Y
InGkLBBoUkN7riZ7OxvfUxz76eRghgwh0CJk7IoHO0uFv4VGS5LBZMM+F0kHgj4w4QM/M5pbCBF8
CvBTEsw2xEr/vIEeLOWpe0nqj3W3ENeOfkmprWf160TiIgYGzBdvn7fxfv/wZ49BkObVrhrg2awz
edgMXX1VsxKk9z4xVZdtRtRsfBstalLnGY01zwfWX7iTY7IRGIVHhDIA4AS7astJFsiFvJvLDmry
goX9TXqOOEV9P4xcm35Z07VBUNeKHmVlRxsi/gT6ZhBjTVspKov+a1jTcRMmqmJVvE4nQ35qQPOE
9m7c7D6+sksE7qP8lugpT83mZuU175IP+Cum/kBwR/ep0WIEjSVq+KQMzM3hdysgb5ELhiyQfSLU
pcu7TFRH5FaUcTQFZssJF1khdExpZq3hd0YzfS7Us7mEbPF/0D99gRjuH7zDysgY7zrHSi2ENITY
l4b6nj7vEmfgXxX4X5T+wUXVWbEHaqAQvJukRY1UxoV+5o8Y8lwptASFLcyxe7MEjoxFHdCpUpPf
em8SZ8drFXZp37NPNvlvTkTjmX3ck3IM+RFMJenZ4sQQUPifXqViH2kjmKF8jI7ELzx22JePxDw/
UxlQjbwbjAiSNepDmwcgMw/mFoUAKRErTv9Tb6Um5xOO9Tc6FQpTn/a3d8Khp2EhIhHtlMmfUOXd
Mu2ORRkKI4lHQEahSd2VjKu11I6DzFYFlGC/lJy7i0CfdX/n8Kjij8kQupsdNxDpRXAy/HNCX/uJ
BoI5FTRr8V6MblB1O7lLVV1bWp6c0zHHwPPFFLdvKZ3N0a6WNygA2PBPCyonfYevMoBnJyUid7Iz
OWTgDeCowucrpN0onqHUq8gS9Lz3kplAE7svU2O+vNR3NSq/Ate2z6UxV4SWODUUo2ZqFrUe2e7a
zDOBI0a/mHoigCBxwGV91Gn6Ed3rzThov1TrTv0gJZxkUGTQsUjzCK47YYTx9+arfCY9fM2A5zGj
+HvmlxFIeZoSI18A9Np27XxqhMaj40uVW9D6y028Pv7k+cDGK+v4lIP6KOn54G/vOz5iSCwDUZfz
Th+v5ZzwDKmiMbqhwdZk/0h4gyMpED49ESv1GBDkJa9wDDtaygTwp5miRFMgN6SMUsc6NQnV19AZ
0d74uVPOL9Ob9ZpzEfBu3kZfqdpfHfS7JFGnhJMwuqncuuv43kqjXOzc5uXc/dKmstOu4bIRvKb5
aD0vt+tYChbBHnOZoXrCfk4R+KTk7jThEOv/q2vt0XG1IR8u6mFc7Utbgj0yUdqasrjl58q1dJ56
TjdWU0JWg2pUVmUTerMLv34x+42K2jZkM33jt7XBjwnVSH2IMneTDOv2TUttQMxmDoaZ3bTXuqpt
1ncaMUEHVxurx1JPQk6gXDAtTsvwMaNikibir4E55yfEUhpdk8kdeItGRS9X/kX0vIKs1yii7TCa
h8k367bXaGFYsAwy6PK0pd2BZQy0ykjJIPZD5z74wJZR6zpqDPIsBWFOp3RYhUP1jy/7dM4SLaky
wkmC08n8MQI87x6DdGrQUR5mvBXFoUkmclFOXnXOWmbnajYMpvgoPSnn5KNMkCDIsBOPT0NaGqQd
ydYAv4NHbtHDET7omMiKKIYjkoDVsDxAaoyABLgI49tZJHOdBGFq9LTvgnhrj+oyAhep/yaeebty
GT8gpZ9jSNkoyiov9QOGWHyn/QyvMjnKOFL3VW1hKaaJnB3iQ/5SooXJhW4t6xREVn/2B45OqCOe
MYzEuwTZOB8+NSDjPM8egLqthaEezcP/u5us6ML4n8lrZhx7LV2dgQL4BvKjHpU6uCgptwlHlEVD
rDjjNUYVytzaKkRQ301MT4O6hPruyaSMGjxXePJkhANAKE08RvO/VXxMPr4q4H2NUjO+ndi1g1Qz
vCFlj7M6IRa+BoGaMbVK5LMmMrWGicYSSinxIcgOt/dpmdq6eq+jIWzPrrVQ2El4eNqzR3MolTQS
5K2YyCdj904rgnY1EHnvGjtHUHdyIZ1a/UeocyfciRNsEQAcdXP1ZQo1rWQNLZMtecorFHyaguko
vGqyoKYv30THD0ouQSxdi17PVVfvFGy8vYln1SDFV8146bMSaigfU0KTQhzrWrPRMsmO2bX4kF8l
nJke/HbHGNKbqgOuflba5Y3m5wAXorznFbCpUSU1OnauJkYVnrtNTGCVlTWbrqcGT3MKfeOtZkK9
bGds+SrNcDu6LNw1igmmVWqnZ87sfcJn+PsWHS9pOVtjKsG7ggoM+CkKB30C9meffL5rEGlHROGX
QSbxR0GOSSAw32czNqHc7nl3M04sqYfY+MVQsobgXyMojcD0+Kag4fJGbEMKzzXBjbrkm3/t38xr
bfRWVtJ5FLvFPJBS6RBSL8op1RIJ8mLl93evNPz++wRtKQ8w5fBwE9hfA9UxxvcuOomm0qty1AIB
RDbCHCyKjeXXUIXX4qsZQeZYsQ9IVdiJ3lDGXEXftJ5FgDgHEtkC0KiewMpVN9Ob1tyNaYACirEv
HnPaAunmueJDACet+0uULtKzwmk1olCPA5u2mAYyHkmWnNyWgZV41k6mUEQcKqYZRXPAffDCWjfi
M9vEtNsfI/gBF4JmpkBE32NOVgEPiKLsLDRQnXC1sv1EFHBfp+g50RvKCm7quo7IZoXfgyzi2jEM
6Pv2sfoP+BbUwidhtg/pFJfiJqIKIYxllPCMHYjcM9CRsSP3TDuvadFyVz1iPcWIgNAxSQ5Lboat
qEVV7EueU8ZsOUWU9oWBSHH4XOn4q3Ms7yQHxLIiOXwrH21C5T0w6uf5LZD6fmeq/z8wqLsPJHaj
3ixkzYIXCbCHGfPtVRS9+ewKypes7KfzFzW7FH4AWM8KoP8rzIp/R7P4qLe/6gHWMAOK/wNs80+m
o6mcMlsIMN3AZbwiQNTKzw6eDuUf8r1jEDVnru3PCwUQIxBOvAE0Y9ilK1cJPAC3uN6V37yq52bS
OQJ6lF+LzeYKbe90P/MJ85svVYEYxny4k2DnPYxEsrzzYwUiNGQtD4+biMJ3jT78hdpjgqLokUyt
sf0Zjfu2/HE/PftyhoiTKCQR94NeGHzYdHdxR7UQHb4bjRy+e75L5e5Azr1TNBvbQ1/LAT/mVYJc
G01slBjCwlSk/fVdiNhOSc9m5401+nrj/i5ybuOpbBubTTSTMjudxbsAUliN8q2bZvcGu0tDKBqd
nnaQQYfjsOfmzYSlHnFDXZFzy1vD2/vKZe2TfzNzeD6B7OBGIQ5Hvq9Ek+YdKJrc1F+whe8U/Gtk
JqX+LP6++oHbFPB+CwOLb50TB75IFLQD0ncErDEYk3RAJ/HklW9Hmfg5LPkOrqS/0I99cvStivIS
FGnhQ+Ump7GgeJO5BfyiInbg+dNTPdNlg12C48QXDP0rPIXRqvbpaZbTtCjIS26O4Y9izSPX6DCu
rcj/6UDP7kQuH4NBGuArYZo+K9WYWbGVGmV+j8MgVUPwY+oggrZmKAVXUkpnK6W0sYYnMVvB5WmW
RSV4FsZZeXhRzAvQX0m23qymeHrHycOksW/h+3FyhgfELjfijas0oduXEAFbP1DdNSQ4whoRyrDw
wH7xr+WyCjAburD1zY4/FygqNGUFjAwhw8Z7DMyfAzpZlYi0rIhW3hlOCBNjiUuZCspXnvYIdeZ2
sm5PuA4l0pvYURjI1BfcGxObe8s6TgLsFGi7T4FBHRCYz3XzOwWhYX0p7V+yt1sVyjpiGfBnomJO
lXWH/lwnI4K5kQxu4foEgZju6+/NGOTyaXH6tQDLkUkby4rx3OwkxpeOicubStSe/i34ZMeQwEE+
co3bN64wQTZvWZSnWHVQl0sZYyKrAZnAuK9hvFzMb2FfmQ+YpmxtQCFqrJsFzO31JDunaSzk3ID1
Yj42RSltOlj8B1tP84qw/TMZsYvK+KubRPN5K0gWJ73qVooqLUSrYwWxzueEZDcdV78Etrz50OgD
5rLLJroYERMe/sDiFIvWnQCM+Hf43XelxATsFK10YCWC1Wn3D2dMJtKO+sjVACt8IkdHz6Bbe4MB
GCxspHqwF0Hzf1CqR4PFDfEucNdI+lvp38G45vepemP9BgsH6DWOKC5KYxFoRe8mVesuc1ioChbN
oK7zDFH3ZEFCZqdZTZHFl8y6h1YYxfiNNHdF4T9mj/TGyAvUJxY3NUfrge5LhC9C1ViEl8xpQKxn
Ay2ls8TaCfYOVFnkiJt5r6Bh0p7uRBSlS5LciC2sLagL408N06K5cE6/6oBdQYkp2TGOz2w6RDtS
ng+V3FUNHwckEyKQs8ozJ7/q5FqWmcGSzGQyMttLlBP7cZaysSWhG8hsBeDM2X3IZGpIy10IQvNA
A/MmEAO9EfCv3P2Eh5Y/IqmLVPoUZBcobxoit1JwRuJl+UFfaP76whU1ZfBUcckHNauHHHbVdX7/
YIYP/1t/qjdn8VxSKhoq5eHxHQ9AcCRF1kjcjsp65SnCEIVdaUeeW7klbXNmGHrgwMXTX1a7NpgL
fAmHblDHc7jLg1CGenfxxANhAFaxogn5WiQ7uXN8xuG6Us0cbK0Wyj+Fpu/I8PIJeGWJiw7fWkNz
YHadptAK7d7VZUXq+3oh+hPMTpTidq7mlajB6VfmxPeXuqWIdOO7jg6UV3GwuAosCE7xlcqWuv07
aX6fnYrG532WhQTU1zOZpVS10PUlU8M5O/vPitKyeEM29+bt0+8Wji6EZtdSW3MbSYvPCzzBZ9HR
AfZWjWVFbVeM+8eXm7gCz2+RYCn0qho9MON5gPOlZDgyp0jkvl8KX2UYJ2cIL6z6uCw6bdtFlTA4
BBORLI240ywk8unPP+AT8uJduZypx52/WBSNklejvKqA8IvPX6VFKPVAv2np+5zryDJcDJWlOsZF
kjD5lLFsDRJzDociXmc3RApfHUnExi8Zjte5w4LwD642OJOKZ0gQXhyI7aWI9sMacNuhedq3XPjp
pmz31k8m6trzosKC0I2fwGWJss0Zu0LbAKmru/xMnMMSwl7y63c6lm1NI1I+7PGCiEKUHTs1Ro6g
Sex0d13Kexir3R2r+U8gDiAI9dgJenc7F33FLhh+z+ha7i888oj7ca+BWf+91RubqijWa3AkdCaA
iMMPuhh1ilxabqIM6yf2UDhIOvzIj2/dE7CEcYy0Yu1vzlvnEnX3O3kIW1i0Ud9Bi30UG7MjcdXu
l0WDIuReHyhGeugr0dgMykhQkklu942ygO9xSip6ttox340y/RvRINy/vOGrXtDxQO7f6AZmupH/
0A5gI+U62Z10tM7IUe48WSM1+uFaCmo7Leg7FuS1c6pFjG6huj/h/3xukWtwmIf3RPW8Yp2DbRi7
nFdeadHTYxB/+ryPPwIXjtzptB/BzVIpvJGSM18aHNDLithY3G7XdkHkaNQOifu0vpqfsg0Vhsi0
lMDSjHdqxMdAe1QV5M2aP8nsCvlo5USiByeJ6G8gQM2XCHNscXifLYQ663iaNan/wFyIY0WwGJV2
EDHTZQmszGNHIil0guu6l7D8ltbonYbJiZLY/12Df+QLpcFqUGmqUWa8iuFTRGEhTUjE/NT0tBLe
Wtec8bAuSG+uGreGFhwFIWC1NYSCiWk63nNWLA1OfyM0Liy63PjYol8MWWrtImtAHRetUC0YGrPN
qy6YTK5Klig17bcJw5AaIuiph9VQ6RTMHm61xDHZ6LWVbhmeEVCB96FebFGv/Jgai4gQdk4Mq3eR
3nU3wCOnPAITJ7s2w6nnXkAYxAcp7GS0cBYjF3L01StctEfAwxwux3FjVuVpeLgjkGIByYtkurim
oO35XYQbLfn5wG366nQGuu3nKQSBLJ8aYqtgeU9W5AZ31OY+5R4U8TLkuHqsnHcHOE9XVhl3+nhE
Id5tqmu+gMfMNClvGpTqTlUYYEoXHENVKmg/FaUbwTqjkHh+Zxm/WwfwDayhXHWtMyqinHoBJGIj
gbkHJtmCFP1tBIRPbjVoeHTY0A6pWSZgi/QzhtS2QOa+5+BWkXf/jec6Xj2eHMz95DmIutSbbmYo
40bOFXn0OaZEVQV6YXh648QmNUtl7LfhW1mvPysPdnuIn2Z3vnUgf4OpefQASa2GUZcRx869QF0t
fQGfnWquA/Bc30ulNutGY7g3wUmaGK3VFHM4AVfv5MfUlOO0JK6uA6DHkqsJVuKfVHZaiRZ3j7bu
7tQPoRt6ObgBOgjKtiwjTNPGIOXZYdniuvwVK2GMElLwgboWfmn5KEZldPBBXXuY/L8V9SznKtM7
tBtSYN/fa6V3Qbs80MBpntSHQMP5r5NNbwAL6pcSqivoMHizHriLIq+lAfGL2WdcqBUCZ4Xz2JAR
bVmLQX89cvZYy6+QBj0IbtllwT/+Gr9LkslS2SWK9Q1aDAVrUY6xCedTaP7RjZTPsNqz/hOqh26w
WOl3Ct0I9uTudd+e6gs6eoOwBvlh+QuIEvV3pDSvwpStTUXgznPFKbyiUGZVDNnLgGJbGsVomR/V
kELtRjx2NJkbaZNdM+T9tRQi6hC+837xWtc04/QHKqzOnHMNqRAcyTFBDH7X5kMrV/GZZ5R6fBM0
5/GYYXfLaSJAGUNoPmVJTfDjYp+iid94DHgLfxp9uPfY71SkCrkK/quuMh1E/6JFBBEnmvfnnU9Y
PDbJGcscfk1xb3hi1waMo+M3xOkuQARxm1oQbbTTcOrIQTSFafKOZADwXhAzvU6sfYDa63XfTWbv
Ccb8q+e7M+6I3AejK1+O1hkug5MTFVa63Ed1H5lUV0HFK1wLZe1HjR6Zb4OTGyk4qOV7ZsqsoMDj
F80mgQaNBTCk/oq5oVawwasI8kikULPBIVMfOdoE5dv10AyIXUVfQ052KhQzGOnV7KEA5JM/ZX3h
5IvE1ThVOjICX0fU6MtoALiV+y46ttcwt8xne9AGYb+VzAH+b49ul3UKwrhFlEloWDqoIt8H1CvY
I0mkJC4vSowDrDXxVTgA/C6wwJTUHR6LDFQGYudbUGaSyjUxNE3DTaA21VK41tJ6CV+iQ6hK/+9v
EgwYBzB8ztkF3ckYnk8fs0Su+xuafl8quthcjTr5m1B8ZSpLrNRveTtfpFIXJiL+ttOu45VrUMZ+
F2VqghNHYU2ry19jfpL7X+b+0Wb3al0kn5NWG/9whiNTjl74rhopqhkFjsXfG2a4RdKSzzybaCuG
e1zPGIBQGGUoJ+u5ZBe5XR7rC7c7SfhSl9PBqa1wIVnPQUOGD0MVYACvZQidhHNK63SycwyNd5Yh
36AnmY7iE4t259TG9CPOVV7MdMWeMdKC0Zk3AKrV6dre6Jffajj1Uze8HkoAoiAl/oN5csMwwrWL
BL5Qzse8V+PAUW1nEy++sMozjr0Mwnozr09JGTG23c2GAgrlhT2XKfoA3kO4ViPjN97fTefHDRw1
ma8euDis0ZijpXG71rmk+XhvSlMUWog7rDzZ0fMy6SS6nV7ITvDxKeE0AOCr7keOVpcWaA5mvkSU
uoWXOCvmzXLu9Am83PW756wNxbs9Rxz7dnwFTO0qIVsiOqj20ai7d3cWPU4nWaOXd5aAagL2W7eY
Zwl6CxD+5FwXcD4S+6GK1hM8Q+ADYPDIrOESJQOUZ0zBVzW9SprVNBHhmJWwpUWCEtleSjhu/Z6y
imkp0J5ZhQlagKbZ0r3tHkIPchlP10GS0ad6oII0hXCgUxr4RjLDJQ+EcjQGWX0bfw+RqQqJLHjC
5JrjVrrbYIc4gPmy0pi1JXlzjDvvWpZPjMJF2i9UB4rwKu4Ah8Td8WA2ESU0E1diUPCNSzPypL70
EnthnpttwzTz+Ju6NEVaEZG6V+2CiKJhGEEuFfZaFbrkbDhfdpnYP4VM5eC8BFaHGsdTXiz0usaC
b88accaw6Ap1VpxtzMBn49ACSAX2yx4sSN4YXP3cEF6WFNZ/cAVHSWxH5H9HLspAvkH8j/i4WMX6
O0hj589USXdJBOkgMpIle73FSCzeAvEr+CA5SZQKUuE9Mc5nKPKgH8gBU+KxwpZGUjmJz8sCJOe4
my8JuNgW39oOAj3TBI5Lwy2KJVUyzIhlMa541PkKaFCot++L/Y7mdVXExmMXoixWdRlWhwPd+JZ4
RO2pOkTIpEyQqDc6yKkXvh30Utpo6vpKiDv5slsL1/hw3oRbIKpXewLoRuzvwwPJrAVyzkH+hQOB
gGJh0cj2BnAh9zWhLqFH5/spwMRFbWHS27OeHxxSK2L5BcnA+trrWO2E7jErzfT+Rz5oqgAudet1
LqrWbPNHfZWNi7fSqMbLVuqWFqj2GQ6vCG9BP+o3N77VcaEY+YdRuGNlcaeyN1SReWatUrFtuvq5
r3BtNQWbR2a6Gaii3LTgTbITIWsHvP5SsRDH3K0fAT9pKaNI7IcJIGgnVIrl0Qn//APPJILME1qK
EyC4tuZJhSfVEKd7hDTMfjyA9xUx4kFjiov9YBX9KETBEKDh4d2gZzi1MDaYTuC9r8J28ukP/jh5
cpeOKuDIm2K/ad+Mrus4BIlx/QAzDGSJxmYHS1rXfHtChawnNj48sMxAkRRiT4/AiAfIoaYK7tl7
pdQBsOI8mM7WEjgPVbpWyBlOvaOFsQIRWTzZ0YRPvABe9bwEkp6wNquH9xEe2VMYZli/AKnaYDkF
h3TBQJnQGYwmTosiFXI3Kt6lvkZtNxMsco8hOAfKoMROUJykdrE8hfXRFDUtqXT0bjOJItCP1Tt+
4AYzgFtUx/K7KbyMqodpkp9t0XqeWwPeYit+m1HQLxsyr0UmgK0hieIW3mai/AIYozcE6aSLk8Fw
eBWNddPb2JAmx3BatyQGWu7Z3JGdiNj6vwL79zMPnvF4OxSrFOTK5TzPtt4pXwauf+4Ejwcy5AVt
d6z1tUJM5P8nhyINRVx1i3ZqXbB7vdgG9RoRzOlOmPn7l6Iru4acIZqfE760t1golMkicvlUtJ3o
ZivwT3EHhJWXNo0c5yJOw4a4821H2fIlSePV/+URtIfp3xl94ZVTfBLxU0GLeXkY50wKXg7n3O7r
QNmdAUMt3qd0+jSTllipcsqYRaLbFYMd8XdTk0WYvN0YIdGM9F2nJ+xjimSBeFTu0WF3c0Ih3eGl
+gYDjhFOwdhaZUfvHwR25XnykxUK8NsSXZM8S5OOD7+7J4J3aWGWP99HejkxlzjaNRTnNHw1jIMS
+VPfa+mlphizVEGKlYwg/BKVZT+Cd2VDU4ZnA93ZDqFAoPNlIJRl3z8YFLZx9QEQN0d9g/dlt/GQ
5JA9Bef/+q/Mj5FsxeVrtf0k4L0aDQfBicya7uJnUuX814ypSqMf/xaTU+NkS6/qn6RgBl/+0r81
kmtmTJMNE7sdpkx/TuB4HMmOsPMP40LkgSim+HuN3sdvLrB3xGhijKp0RsyFMO0XhVjMTygslJBi
rx15qob39hH81V8cwosXAbTzzem9LjiYo9MN3mPdmnDDVbxKEDWsid5LPZ2X4PTeKRE5wPBSUsSp
zZ9gV0yqjZJCBmf1ulEEtshoKWRU2dkCpYJAhw/PtvJo2oy1UPF5y0urD4TOQgPrz1t75eF9Fh1t
SHatf5cNIdXReJJ+u3Nmj2NOWUto9n0qEF5yHeDzEsQ0S1gTt7MSAlt2ExD8qFPn7gmC3C6QMhJJ
/KPhh+neNT/2REz6paZac+LjIlmURraF79u1icidBHIO1Nxgrd2VzDed+oDWuDAg37ig0ODQaYkj
jhh7vUQlPghNiohruVuJuw7P6L0mMtaaSQHb4zCpCAllD8gMdx8bF68ku5IFVsaaOF8oLvBoUR2G
9jVinBJuR1Wr/iZDqPogmg1mebZaLy7NKOUWs1GIH8aw5G4Y4jOgoVzXXPM8KG6sd+PEkavjgUMJ
0/u46EskDc5sD8C2odARWHFCcXokRk8G+6YVP2NqEwHGi/Qg0aDARqoBkwEi7sn+Sr5/9tk62FQ/
VPyJsqX8uFFX1BXJYFlGa2E6IZxcOCt/TdbPecauWS2fXjFJFrCx7LgxOJ1r/xq/ut/bew73F5Xc
ShuiQ/fAAtstayICUgNS8sog+93jxeVCBUXi3h8XMxzOtG5I4lM7oQ/YfX3D/1g9G4ceZarezGlE
Bt7EGuGmEfc+YQueG81LNI6eIquMeGtkM798/K7R6W0qlyi8hORt2ychv4+FJFSXl/eb5dpQHI8D
6cV+EynDnMzRERJJF7mnJV8eCE8lkXZ4NMDZIjs/3fvqoTrr7EE2Rxwi3sYtufSPr/T/TMnzQpSO
s+UDEzzV7HWPDUrsbzfvGFVz7rte0vFj3gSlo3EiKsrlYnbXFymM/YYsHn5/Gsw8nf9XzHFiD3HM
TgK2vEJzZQn4YEyjYXGoBR3ZIU35IPNsPBa5RKviVF167Jd47sjIFh7WEGX9EITid3T+jNRQuKcn
gBzUl2xOuKCDqtVnjQ6KCtshZ/f9s4f8tINNd2UavhFlCCqIRiO9glJOIoOQ52onGSCOIRiIz3Gu
VlRquQqjbiT/b75Rgc2ZbDRrdQqQYx8c0BCbTU6Z0ijWjTd4/p0u6K1nn4itinM3jcNLpHCxD1FL
Ne2g0132Wr5VJ4Z7NUzzVHxMYqePZeQNDLkQ9AG4XrxCMG8fLjuFBDY2c8oVBWgaSWb92ioau1sT
gzjAQkdmUCRTJh3mv1wG8DpmIN/ZI+CCR7nzTgo/ikqdNYJ9t0TayfYsUgsA56ZvVB9HllwhrWRD
z1grPy/tawTqEg++Wka7Ie9EBCFpqhFiWoiR6x2jHHgLXrvpYNYZlMB1NnVttHYR+FBEkCw8u+5h
x7u9gwIz6IHwZHDAQFuZ9XDqaa1QrInpfF+EmO7KL21fY1tRIf7AWzoPBobCcUqYwxO/C06IuKir
PZaqiT5E1I/NGCivyzRLVo6w4liBhb9sBwq9+zHMk4CXHxzUY9Udlvd7J1eLbA5eHRcN76JYj3rk
T2WRurvMLhebJN8NzTdGzSwneopa3YRDbqlTyuOcX9iDyx4TSs5y5CtTF2HtmiIyp2lsxCtXHvI5
LDRxlsxkJrH8Lk1ydXOKt7oqk7xXlJGsGEhiqhNGOxmAbhizXDjtAB77ZDRopufj8dCFZVWaY0ua
W4G9jITzc1GR/n1HyOqr7+yQnrdbdMgKXGFwU6WNGC1wf61YPjQHP1CBopGzlTV5uyTxN0nyc3Gz
PsfRHwc3zvPQA9FrlY7Ovhc9wmW+dc32p5p+pBqTh0LG96rM8HFbDf1p7le3Xpi2aScQcQA0qEtW
7tGgYT/9Krf7DCdXvBjFD2kxNEDG4zUBJfm6xvgBesxqOAOkv17kGKVAqcjy8A3gakT2gy1XgTP0
YwpxMxsxjPtjmh7eWe4S7eHyA15d+KVZMxZeUT+wdHfYarsMfYToOtslgUM10DxE2Yf/4DL5pYwK
fUmpjKA8mN6P4YZHRMuLA+EZ4rfWmVeCsMq2njA0lDXBEybIEFm9bwt3A0/Oo26/qP/3cNFlDVsW
I5QgnZc52xZFy/Z74gzS618jHtEl/kVrvmdRfgIilgvr3BlGJ2iJiqtvOzlWjiJctoE8lcqztB+A
DSCAng6K0XpWu0PBnhGTHHNqVi+z0jKPOigag1KYJDfZQt0fdl7pnVH5C8Za8iEz6hvplazJkOnh
sjO4JtyXv9avJ0ZAqrmS/OU+nrQ6p+uTblYh5pjAysZq7HC55jAmHznavOlN8WRoCbq6j2YJoFAn
Nz3n0cEeWcneIpu/UAe/U+JeU//qGEzGyyZcePGLw+s9bwCkur1YFnlog7SwNd1/UdZbwwACogez
Vyj6VQShQ+HEcE6JY5+4xuk/q2o2BbfTvv/tAcRkrs+qxOPI+TQwxZQHe8lQ9uc353fFdsttoGUs
s+Il1kkKY+Y+eK9snr3gIydtFZjp85gWlR1lqe/SkvRGkBnms9H55odvav6ODGgeKORAQvbJrkn6
ydgta5kKBf9PlC4AQXEWwkto8LzbA20=
`pragma protect end_protected
