`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
IfjuVOxx0E7myNYeV5vc5Nr9aUTdgJjPP/w5FyNj7+3nGzAlGeBsSjsj18hUaHu7b/c4WtSxkgys
0ZehmIZpRg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
kyCZJNqKZYiw+if5fQQWJaAQV6y939PWIVdYzhlkhpK/wIKRnr65kteUauaJUfQu2nF9idqt6JGY
kD0Z6wxRORZicW9jlC8wrCYdslx/ZdVfOv8cRZ18SPY522/rsXMxyTuSGU/tW0Ca9fRkYa7+BCWj
jGlsveQDkflESVcRcNg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
z7LaeD2O04f6MLEgRYbSilNz4NmoJ/R59OUl9IN9P5+RHUNw21MzKaj26S+Ru+785JEAPBB7rdqD
FQB998wBvNTE+QMtEKqsJMDnb7j3njOtWsKc4f48nitm587ZhfsKnajWll5f3uSCpD6XhUrgnrHk
iifpWnfZbLZJveectkhnYvEcaaM3kIuHb6thFb1aTjqLb2P10jthyVucFK7qLyH+xySH7YQ5IWGp
oykItTDPEFBGo20Wh01Sn24cFCe/8sg45cjFbREqqNy9Aqu5/DdTDFIi7Dn/LHUvphhtYtVAXNzC
4CbAI/JV19rthAZlDEQFJiWBCZOtjnOO94GgNg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
c80d6NhaoF0Fw2KSX56mwPFk71g3lQ5boh92tADB9KbWJ+W3pCXYgONMjfElJ3qxA+zB1dTK/wl+
DtGAToJKTVZHXf8wvTZxpob/x0MAkpvwMKSuRGUa88ZL9INFp40rBgS3ZJ1JeWUPtpLCwNWifm8r
vwGkpkFjFpU6Vwya0mL5lNeJpbc/xEFi486ohcm0va8D6PSk4bjBD7o3lzd8exDM0hbFbxZshqDo
NbA22NyjGv6/Md1D1Mlz74o44biX8SzFkwBLk2uMAgwIEG+suA600mpOQ7tPU81jD8QSRaaMlgAO
CNd9elRv085IoE9qR2Ks1MkacV8ZYBrkNbp4dA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
raCERu0awtcm5u22iyLt0o2w3wIsu+WzGRUPdEWE78PFHKGYcEx74i90JHjoo7REZxcfGnyEXPJZ
JGVYZl8bj3AwjIj2hwMdUXApo2y7/DJNDWdPLrDpS5XWocULxzXN++C+MWcz0p0OFxds46OfIcY8
abMUKhNtOAtyRdd8Qi1oIRJgyYoHuRwu+Vhw7xxLgVrTCPFt/lP+b8sQxbD+WBFoSquQRJKih11v
Pkb4s9qGoTopeqLuVZvRm+CVJkXLrZaRaPPBoPVpv6H88t0el9WUJj6gKPsyxop1hhCIKuXJBH4F
7d9F0pc6juTzI9W0JE4M4Kw3HPBsTDh3UInlzw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IIdGziZWkSTRRHnODVkoEkOMqdD2D1/bvr4uVbRHLxk+gzFdi/Z0iCVSC10XTpbZvt5P0zzLdXBG
+91DTd4vXkFBEq75gshG7o0Uekci2HOTokjZQValdLUIJJGOfRXnYmYRBJtXcSPci8llirCsVqof
9Osu8/h4QmeLG6DyylA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FlgxLsgJw2fPnsKtY2d/BZIeMAU6WZ2xfe/3w7gSX/jJaZmDRqyxqczwQiudFCeHF5OR5L9Qec8d
u8V8eU9Upe7vSl5ZNFEUVqlgjrNc/Y7OKNrzzKY4iSKNxVlV5sfO5YwCdFgq5aUEz/2OX0ETEmOS
1XTfdWTaT0C/LUwtLSJVRyhUCCXahQ+aocamo57fwknsXoWbI/UbldJi8ILttwmQCiGGTKdpv2jk
FS8mpW4OFbymMBQp6j2JvPeJ4qRvFz8X0U3h6sPXc0bc+8mr51E/O3DoNju2Eao/ysVxdM6WQyhQ
5HR6ddheC3re6Y0NENqzH/jkA3YMv5fjFQ/DLQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
8JsIwqAUF3c9IdmDQRcbsZa10Ihm6sLPxvyOm0Vl/yoMY01TNhmPMu0RDapZqtkYghSFz9DiZ8IQ
rIme0GN7xuIo0hdidF25ogTHNw+Jb/iParLz1RfjOIA8QX880/goL+8KKVVUOmHz1vQxe4sl4SPw
cJO+fd7LsONpqxG3MaffiZQcDpHwD0hcijwGoV2x5ZVXn2VYnY3DHIu5nqjAvLMeRyhTaUo+Muu7
l93ixYrSTWS3Lr/7JmP1LkTPGLziX5YhElAmSIS8vfCtDSKQlHLnnALRXTHtGpH5IU5NJUgNdr3F
gJIoxS9LUNJhqs5VaIEY9Ulvwgiwq3noQ8ZTgUkPUKM8C0DNf6AVd67xqyrdO4fhUK/EbFw9G5tH
y0vTzoSgfvoA6GQqEvk+ryHc6O9jFmxJOWwK46s0IU8yx5eZjwq8/wZ7Su/Px8Jc4VLt7eAhKqxL
rO0DFqyhKUr8jhTt5zo0RegP38ffW6w8ASP5bRGHFHU1lcURysmznZlTXtEc0u6FCiMA0x5GdlfE
zep/JyB6BK2f7ofV+HuiUcz0tjkkiKKXIEk/9/ucPc9MTL1MKLpAkcY0waEsD81jcTuKipYZQxXJ
GH4Jnk97ThL0MaX3EEut7+MDjpMrczJ7GHy8eDIEVbF/EtvM3mmp1qRHewHVbfFlPCH1qXtb1NiU
tZeqNqwM5dmiTGD3Tc5gn/gyYJCwMewEx1NNAanVaFLe0K3Izb09bxjrqvTi0aSywVqRZXK48gDM
633WHtjDDqjnDPKKgYzQZ6wfZq3OJN0K40ZdsAdKq+n/L7LanXVDxskAOBw3RNkA/EA4IKzLbp74
izGahe04XN5KwWZLECZLIoFqzlnOhc9CEXYxpa0ih9bpZqsGhQ2jvM9v4WW7EhnV/sVI/vTMv9SY
XBI5AdIrhY2wA2R5wZoZu19ylc5OPV9fJoi2R8m/4O2i4y+oFcxsJvAptsCCVDeryewy3+wX9me+
ijhUv0XKPzlnrHP+S2+AEbsoPJWBhJkqoE+d1MTjmOLVKb0/moxFC5a1nAb1Cgs0i/G2H+rfYS0f
gNp4C6xlU31wBN7AyCVdj9wl/lAv8/dp400VrNRYnlr2HFoDNtJBqqvrOv00yGTtnWeZbgviwY10
jIf2sxmS4uLuehMlETDsInRnvz9R7TV9iWyTEzMfGVSnKqk31RTlw0yEoJy7Gt8PweGDP/W7hX6Y
9Q2FOFmxaQ8Xp2CXQlhvnIijIKXiJiF3+T4SivLq6ypdnGEHB4c8BV2DX+OUvlD60PsVy03u+C/o
eaqioNqXsvTIzLZxbxsdkBa8PMzcv4prZlYds4ZrNqBKR3Gt+WOsHQabqyQ/FOBfLEjYtvDHHYvU
sq8hVj4ve/3d3iT4owO/5/ZLKA2SWc4gYF4mY2ndIRGVPYXjkwZkwrgxokEIF+2wOVA5ShceHTzv
SV1nhA3GcsoN+VYfau7SDqFVnGh/nbZWEoFw2H93fKMNSbZbsO4UyX8S8l6UT+mJl+sGmZgRcm2a
YgKr/kDNMZpuTJSK4nAbR3Mjxy3wrPlJZne+UI4rOP/7D+uvh/aB2Du5TxoVMOI3RR1EOKBTvM2k
O51IbDwJLk2zefmspKqGnnquHnsTsLsOBl0twtg0xxG+TYMj6dk7ELGz4t6FHZHEu/a+Hdqp2LX8
knfXjehiMhATPrJ4UjOVvoGrJ30bvKLDVGjDzJN0KF0g7Vd0c4i/KM/yOAa+VFE7VyiglU3TbR8Y
SQiWCHWdISH53339zJ0D6WxsZhKAhyFMNBU9RgnxVDDqYZU1fGJoG98QR/kmcIiOul0kvrpTZRoW
qv/NYqN7O3g84xO1dUyJvmXHMRpbl3i0rhehBeBVGXOIpr+TNvCHStZQlorVFKSm+186UTHb4UB4
ar6iFkUDaNuG/+U2BXfV8mtVDUCvL79RHvd/LZe90dVX/x9RtxTlYZRiKykARFMcXwXnZeLzBfqC
+PeK7r+zafFTVYECZ0b4UiY1Zy7fEWyHchETe+xJvOVGajzb9slICiIBFx4yc8IQyoe2tenAjqbo
eOFGiHz/A6PbkS++BjWH5B1+2HZg+0c7bE4yfrZZ67YGqKZaZkOKXY3POjlF1p7bpAHaGgwhyRqy
KJZuXjq1QXPLVkhgx0vrCKGz8ywpxq0/g7Kit+6lmnnNxgRmAd7Nw7aLcIkmMxmB778ac0WotAzv
QQ/2tYdU2o3XBSR5/ExQcA5te0bHSQTIvWJ/vKVejRoRAFi6CvhW2ET+y9YJS9DOQ+NTQI1ZGzVn
2dnDuErhJoX0CE34veeMT8vP/W2mgJyz6Rke9JV8b0k3PtXRMN/PBgxM24a7KbNyGYygUmwpz54t
FLhkP8v51ghh4LMb8uDpC0zh4iVlwDpYkScvsMOW+uZfEPCi1C0aBZhiPi+gGzxOqNcBitYdfM7t
tGGQjr1P1Lo49R7FYcE8uxHqwQhGS0R8VXf0s9g61Bqr/atp/5iLq3djqjk5xPtGNWrOuqPZnaRj
hPif0Xd39lJRQoNdH/bqIVN3/7Sc+CjIzJu4TJc0IbQdiEqaNBCElcgQVwOP758xz6gw2+sBbi3n
tpXNEgmSeKS6pWIvzjVIdsE9MQUTiogpxXh6lubor0G77NC19Hx/khP0uMunhb17qWntAXY9Pj9y
rG+TioDgXsqlgAttcuvoGJ2Uw9N/ymNdkiloMj0l6JAOhLyxzcHL4ARHQGn8Y6Jc/C0IHbNxeL3v
dC4f0cY4zbz6Mx9DRRVElIvyraODYMx5gsDzCiQKClWMFQQRRZYtJLSXIH46PunSDpQwe6dJXElN
V/MeSaMWt5Rr08wZ8u5hBzCi/t5KXsiRvtAgVIhPH6auwlcWYgtTc+cudVn+fhsGIm5yDyijr8M1
cYLoLFEVbv40lxh4MsEyaBileZvERVCOKmqe9JR/yjn8VIWOt20rQ+51BOAbURsbtMBF7p9dDAo2
9Dj/QXM7Qe+AzqDBxSZd2o17aI2xX0it4BQIbMwCx+ZrNbO0Vb9l/YkFx8XD5d3IyyG2hk5zFi9Y
LCOMRznSlEAwJQnUaypb0mdehQ8GXppRdeR5fodlzXjUheklqE9vGZUyfMeuMYrpk57Yc9NBhf1u
wVo3QodyByQqk9AV78CHwmojr0JgSPgY0HpGrYrzjlG/lzmb/Ozx9I8HB5Q94mV4bR9rneSurB/w
KWoyECj5bk4z63Rh24PHsDYvlHxM5gn0COZ+QfYGLd7VXckfNJ/VI1P73jGWRV8xHipzGzG3HciO
+LIb/X0FwWGy6wchYIKzVo2FuTb6CK3fDiUt+ghV8ttAfamPZXZN4potrG1P0ZZku3wLxILhfKqD
Zd5U7td1MnmYqHtoyPR5kvksLupGe1XDEyBsGEZTkRszz6MBoWmNHmhe1p+4H3TZrD4F1wBmZy2Y
Mq2VxQWhCnFkFYHwZSZ9WWKGR+LdGCZLe1JW0pUSL0O7BmtBYRzIzGuLxJfTOq0XFjwwMseQWvxr
kvGAcOkvZ215kga/GiKhG1CoA1g7bs9kg/SFKa2ZLjRypfnma2G7ePKbuaudTQ4T0YKEPbJfjFkR
a2EOl8jUSQPx+ddI6C8yT7BnjmUYufmJwEpCkm6+RdJzd7Cytz2rolELZqqbwQBtk35z/PvfYQdg
LztciOAytgP2y5lVdlqatlUrp1rwWZqvp9TgEt7ztMPwN8LbuszxVVZQ0Thw6JuKYcb8n+EyYfOd
vTwPuAM/ICnZrgJ46Ign4/TL9H+Gl+CmIsRNI20Sx11chQrJ4Zq44IAIOJiDKZhVzRuvsJKOX/AJ
tlOdMsUD7sMUnC93+4P5EY7xpfHh0142Ps/znnPSGyU8Cpjk1cta1tpaZ9GA7wYlVbPmFd4lCTyb
wM7G4GPf93fhSAaKnOB5JT4KwlPR8YJ+2UZrh7SU9CVFCc04VIt2e7Qx6Hc+U6s/vi41t28ECUNA
yhUH1sL9kaTvJg7pLKUE08kbROoszJ8nvsU51U/2OyYxzGw0JEnJgvEtPunDDTfAmRhMck6YCfWb
wYMdQcvcsI7lrUH1baWzvawHonry+xK7e/mHKLKY1GRlQEo6ahy/IsijukncDGG5IqFCMByGJVQG
xj6dJUHudPWmdXDLqi1cJjlCqHbSf5IyN/XLk/3IjdCxOvVqQGim4wUpFW/9rV37QhJ8tbQaUCC/
DxiwmdgNITHA8fxRi6IiarI12PFNCTe3RvrzRcL2m47fA7SgfBOwEi+pcuEkvOUHk5hDPkajkO38
iGuwKIFEeJZccPRIXEFqL2fjmt26P7NeocmZ16Wkw3J5h+Zvm871Is5mQ52jI5YGk9hKfGfnfQSI
gOLMKwVwaqapvgD6CM6SW+QbE9VXsd4SnQ5fUR6yyQoXX64HIt7cEhwurblL9mqkZcXqnDCELBCE
uKISdhfPb9EHGONr+CGV5ZbAJsFOYy5hWz7mnP65XC591XYUXMelskEpo2p150i4aZ0EeLFejX9t
dsaeT/Kx3xIdctYqwjh0HqRuIr7QgDrWrWX6XT0OUL9nJsUJDTVdHYRqUe47FZlmzHrYTmPapMXX
oUfkEWgd8k9I77J75sub/W8iC7o+RGSNZW5qdJjOn0vKbjhlaCJq6ADGR7VW93rdEXkxpciFsRFp
yFI9LYuRVJasJwXeg0wHWpBy7plgXrFG7kWR0kEy+h6rDhNGLOZufArmIJlkRqjr+qI0PwDbSHoN
mYYFUpvVR5Dzx9+ZzQdphyKNpzcGwQwtzZv60StHTa9dJf+fH3euChNzyB11YqvR+EPnrdgFf3oH
nluhhePay+76EEjICAKILVxzLtioNdOxwC6kPwZbmN2eeDzyIjpcyv6wZhpBwlOaJL+SwvkbMcrW
349lT4IpvvaRLnJhrCaZ+GA3MR4wuaMWyW9CzX7v7EMk2Pj273LZyeEk9z530ajd7ihIOM78U5qv
usSR5ejaWLDerinIWqshIprb2TmrgIc2yKcZoj4x5IIbtX0QrDun3ox0y/B59Dh5woggUSr2hCA7
GGLVZGTSFddTUBIBbKSRMDOkQkp5GLpNuvRbqYXRNqkFK3pupRbSY9XJBQEav/KWrSrf2haE5hpI
k+BUM2JDnkXO+xTFQiL1QNmwTe7WZa3rYtSzFejp0czmacuV3+BGYETCsCphkl3qFKKyyLdGQ48l
587cCzP2N9pIxrjDZjqcz/TwsFPgDv9lQSZOQBNNdoJeRyhXGfGJefkE/lmuC1qvESjQi0v8iZvm
VZvmhydjpCe04iPwRtPB/OlUCWvRodusDBFa+AAlqFIqfDjyhxsguNHReDP0cO5qFGfw4dKTO6LR
sbjCS44MO7NSl6TTM8360IuMJH2H/fGawjrffuIkPi4vbYhe/ro74O1KFQlPbUivjYkoQZSDaOf8
v7mRpyuMvyZmw0tXZL8md3mUNWdT+kesbG1TNgHJzDs7XzzbKxlYGBGf8hc0Q0VfMxyjmrNcnAKe
4RjorE4nDx8yvil4NdhwIB8lK19BkoAancAnsydCGtQSd8vZslcmUgdxLZr7HFQNgYKdfmb5GdIF
FOGD0HVTeuQ83n6kf9Aqb9DL9NSBhEnrykz7k7VSFIQl/rxwbNLXwmZ+Kdd9IWHpkniyybJoc4pA
76DiSSQ3pqQYO5I46O4CMdD0rzI643ClKuC88rR8PMt3mNBPxeI+futs7uwtyvXSah8B7mvK5ptb
VsReNIFx09WFSbksDhff5rEzNHOOgp8oQbn5G4AXuID2Hrt4Q+CMHkZ6PmgHISf7qST8tYH2eNI3
VifejK03bvWlUSxH9pJ83kD3nVGH1PjA0v1wRqQ8tE9WSHORzMsKbVq6Py3cEuwqf8dDSjW3+3QL
kumNRL/Cg/I4OLS7sI+HkfooodB5ThTdWGqNC0j5msnk62yRm9SQxT+JyyNmJBl1AVPe0EbJI+0R
GB+HgiTnBvhYfc6F5jVKEUCNUybUkis6GSL5TPTAB6mRY5RCPmZAfKsqKA0i2YnDTzrTUaazmnrw
uzi1P5J4uSWS7uWiuT2hHaGKU+i9OfT2jz1/JRrzUJb5HaS3EW5mZwKEOKllooCeuwqCJwOvxmTm
cV5OXyJgVI3L/DAWFbvU+YWyuvsooRqWCWCBhWhUEEDyByD5XflSd3v97Yz2xg8eg1vVV5h+hVRq
Rj95AVoLkcSPdlA2FgCaE8Mh5GwR3b/urcCoU1c7chxB4Q8b/+nocZdyriHh1RW6uktNpaajNHGp
K8ufZnEY+qT/1OoL462q7iXVwtGwJHI1RNrJguqdnEa/SLuwZxTQEGd499Nf6OgPisSEZkghIz3z
Io3zznfjK3V6/HVsfkI4I47gQT2yCNnw/6lGPx01ijczNWctoQmy0AfCxdj4l2FhOitU8aPDq9iv
KGmZqOKefoyn4VjCAU6VBoS/a0pxUmXup0cgRynUhXL955S3mnD9rao8y4jtFaFBPUZ3IoxbbZys
XsYsDgVr7C7zSsBYqv0/4CI9ths9Wz03GNQmIBPhKFiCocXNwyAQ8kFZvLaF8CvaGnMwm5CwK2h/
SdODEKTcyvulmY4tGLwf/iKa1XqyxFQ7/uCeIVcC+beGSc7rTy8N9eTqzjRxXl4KgZ4UU7p9meGo
mLl4gigxdbZMc+P7np4cJhxgIFQQUGgbXFsBXCCS9bWLzvYFlQG5XNS0bDmLwRLl9GZl10fiR9ND
Qa6mmUs+hZA1/ayJjIdpo5zsU01FvDdLVSGnSKyEOQ9OskngcO5iO2zCpGoQOeRvewPKd6RmfkrS
Evq323PBvtjG+5DUXa3Dls9xLK9bp3N9ifI+egvYwAxXBqvo+rkZvA2vTV4FyOLqXoxCy38YSSIX
2pNE/Fnoiz0+ifecy3swQ2+7qKqMBmos3zuToPJ7sv3UnrJWP3gxcc+FaP0imPRONyvncr+McRuA
HZuIAvPjq4zYfemvAYcNh3+jvQk4HRAMHTUHlt8+l13csDysIouUNA2iY0iPcFGMsUlZxw7OAwhg
iQYAii6LJRutJ8p5aXP+dXGSJpOuoFGAhgyCaasdsP0+O+Qob1+W0swPhNorBeZj9L/dM+MliJe8
JNlzv4PLJkKsMEbglvQY9pUtkLEzHLTBIeUTFWWbEWhZdXvZa1mTFU6xKVkxgGWWtdLAzdoB7Xs7
cPslkcnyWCHvFbJeZ21CYSFTp7v5eI7W8FT4orbpQKijKHe1YLbLCZAXYro8+mTS1AMAOjcr4JHu
jVTrKW7IW+b/jntrz1CVK/9fO6gnwnYhRUexegBTJBf6SXAUNO9H1nBHVLhSo+sYqy+MryWNq/8k
mwp8ryNXUWaEuCe91b76xADuE2dVXXJsKmvlXXnd2qOcDenGY/noJQRb4/Rg4k/8xvQfHK9lUtyY
jMDDE6auCQ1A1nXjVUZd5ssowITH/uSBHn5dudUYtJ8JVbIV1c4y5GyvaOFpEf0w3i3I4HcW/FLM
NnaC1Fgxtr9d6jwSO1YmmSY7n7w/7m+83PVkJ4g+GQGR/ST9SlgG9z2wdVNukqIdQPDB9/eodSUs
VTk+GlpL/+FdAMkwu5Gb0QckNuYCwFxIti4NJ0QNibdR3we6tCOUUaQHx0/fHoKaxhEwJTIhtIFP
tIVQQESr+nztylayagnlnNBjhSkw2+c/PURwPzoxns4PaGDadfFGI1hYzhFzkkldxISa7kOJjxW/
8niRrNs+igL6ZzHYSLsHCg8fySc8tyH88/l4aCCtHLJizcQvGkGbxvkMQmeHjF7fOa69VcNtV7tZ
UpQxZM+59kS1D/6QV6aiMOu0FWT9PqInMdyKjbc9ib+AF+/pSFT2RUpeurI2lNb2dtcM6a5Oo5JY
Pl7i94PoDYyEJHMC+ICKoTmI23RWUhhQcxyU2DkCl+3/ta12zxzOBeAIj/dvyh6LfnTagzH55Yvp
B6icl9QnaKxSQ0XOwyL7aPXYfiBbk2QAbgzSv2MrpHsdbbQiOdcnCr0sY0c9FNrQKseEajeLVrme
ZosMvJ8CWt2ZQ8OWLuJ3m6hU1P5Gnw5vY0vIl0TuIUe9XlPDK0uq33uq7alCrYiLhb+UmyQAr88M
tsXlYP4dx8HG2ezpGc5KYGbE5218O2MFboXHvLOvXx506Oj1L1hDOoD1cLMJ9Jh79qQZ63INFoz5
7q5y37llm0ziKpJTzD6BoCJkTb+7ZzX/MRB7HQFLgdHpVy6Y/MCs25jOUUFcZeRpWtuCxD3Rwumr
QhSnRtxtGyjJXO6ua+gybNDYLJ+i4n0ugd8phZbIWAW7gQywCXCp63tVd85pkD7gXFp8+SzmRkDD
g4T5qWk86fO8T4jm8xL87r0ZUubsClPN3e/sVVyGMc3i7yd4G7bBcm6AeRH2CHw7e7HMjEG+kP0r
KHfKCXyHAYoS9ddq4glpo5PPnCqTaenX27lA1rAxElNicaVCvT+AUk0vnNJQZ/w3qbEPT5f4Uoo8
xzC8tqCPxpA2vqbpuTcHNe4giSNI63HyVCkbAi+4bQ9bWws9FnuCrtmP2A29P3QvyFM4ZlzSoDP5
O26+ropK32hmtqaW2In3zY7FVB1bZhbBRDcOpOIizi5b77OukUwTxd6YTeAvoLsD3Rl3OABxkmbs
dKZ8u27FggMDtZb/lE/KiQw+v7W3ha1dnv8/0WSK4zKGel/pBsr3j4ZpcJB/7dbcD8fXOEuas4ew
cqd0KlfCQaDCyMiKw3vBQ+0Tcsis0J6qWtZO0/NJJ6EcjyhbEI+WoNqBYusgl6kNpAZHtCYK3HWr
8gWF90k7CzPk4sCwJUxy4vh+a3kLKPcFld0JTer+qEWymFlxgKjK3nr3EmbuVUxazZQ+bvkRihM0
Fjte8IR+FL2OwkKN9BuvzBgpkXnfK+zqSXPs59bFGibCaIdAE1jXafys7At5TGu8mYIHqKp1ggPi
PZppBZJ0qNmUKywIcbO7LImSjZFfBuFdD+XZAVtdBdB2PqYG7tBEU4EbzMHkRX7DcHW2wftw8L8u
cwyAFNzpqJw8IMLRb11l/C/0FGPitZEg4rKFehLFnQw9flte8RWdlmY6vxdwkWd3aq0SouT3V7aR
mZNPbraZ9c4Ne/yplDRz8+MLP1RsDn09VksPYHv9B1nB6E49gc66vrIpQce/B+diMxvtgIbTbwhS
G+EHzlZ0wMA21MtNToc9OvLNQVLF3XR9+uXWXF+uYIyUzCKbUPVxeqtTLvLNhJEg4wEcw/JXJYpZ
M+pIA4NlATOg1uYqTivRHOE0BG05a8/Y771h9pqTrvpop2cdyVIxV2Zg93krRk7CRuijY9334Uhy
UYHnGZjgK4xxnz6/WHj+/+eICP1Q28IVthFishBeZ8Ir1nzBvv03zF2NpaT23TPTRZWQSIzJmEjv
SXEsTbRPnXgMOLgjwdpZZnUaCIEs1QAOn01bJ4AbCOH71KzFmMyli3ewtc4lrLHKAsjLCRrPfO8k
TT4qXwsTwtLtjKQnA2nWPQ8kaowVpTHkDgm+06/Zzxp0qxzrbxxShIyp4mpZYziH0K4dl6cMBVoZ
C3uCyHt+lZggS8gZhsJJZ2AitRethn1PEoHVBKNPWw4ZOuWyhRa4Gk4H5J4Fzox5qF8s9NBPWgfE
CVfnzPCQa0k1g5T1B2K+sRSpaBVqXPcukHLA0fBcoJP/2kB0dKpYfbBfLz3+G1R8KLfC7yatSyHL
Qv14ECK+VOPBcE2OPtBNkIude6eOZw4KU5dOJEljJgDqq1ia53kym7xwQiPpFr+1DUxJNfLrz+Q5
r+e4SC0u2BaKLp3hleakTxZHQ0nUNSX/IX964UsJZdGPRyXVXbgSDQo9MHIGzsV1V8bpJbkIJfGu
f1iFkBbl9KXrfRcd/wmstyz+iehcwZeedG8jRIzQAL8W92T87HJWwZM0kR0VAKumgNRju7ZHTahW
vSJXvlh8zv+tuHRCrQAtW7Kh/jXEJ2pEMvzWO7PgaptsXptP3MWboLwizqJ3n+2hnmlAR+UU25oL
WNNxdThnittr/XXY7BfQtz+XRhT0MxfQb92+tGjDTkzCODVX5zvjv4gj1rmESt0W+QjfqfBOubas
SsViW2ltdOCZ8QJZlw/CAFCp+hOsStR13iL3tNVcMMKgpyqaaKWpMxO0pWgbacrDNT6iOxOaXh4b
BtoGcpaDqp+pDPJ6QBcEFvL0h8i1o7uXxL5b1B5EZWPul7RcnnoKyn/qAOjhwgQKuIleUa3QMgq3
gB207uJ1KHcl+y/Ygy8H6v+Kd9JIF6J1Tsp5zG0yhAKDWpntiWYQJTOnukGHnyAi94tCbekazkh2
omU8B2BlvhMh8DbJHA33+licfnunMbyzZ+6Vq9cGHUUP/4eWyJfiyVc4436PeFb3OkojOxy4zTUE
aro2sbgRCr4lp7RpcycQFjZdlPrYRqUnQi6OSUrNgApiRNmewHycWCM0/9yp3afwFkYVRoYp/a2A
zyPlddfZ3wNm7sswnieXcyvStaT0PstAAcxCL5OkTCWF6aJHAiN9tEDIccTDeeuCJcZFYO+AOEki
gbZZa+LkP+pS4OV7PnYLa8e2mhygGY9PiU3URLJVGmZwmpuVmDf4aCy8Eu9AOB0yLfl1fKo5/vFU
jfkPQLFl9NzAvr1xS7HSyW8pqPEAd6Kl+NuytwxlZPpJRRfW1SGJ0RIuw9OFbxlsgt4A/Vjwqx1P
rHrePJYx2smIbyqL6HnxlYKdAwyQ6h1a7C9vtg8I1XMpQaz9tlvlaJu7BXnkU5r9oQkAxBiisNrV
IkhIq55ocvPyN0GZjIJXxQhj0I3hNaBv9ZL6VKGMa+vPx3+O9HAfCAGmbMBqFamI2Rj+0/AEsA3g
zsOzgDMzNMMfmgiFIV4C6YiQQD1pIv7SYVVKvVoVbguZkdGETFgXLnIsTs98GCMii2m7mbcRXh29
YqGg1l5vrMwy+WkxUvrnTICfRMRkg3axj/A9/D1PJbmug5PDT29NPxbbyT9IxJt6Y+zbmrnxLE4o
ZC1LieF0Tc+nC9c7Lwb3zjltd/3x1wTDTq1Lp94+4Qk1OY+DAn7KrbZx9A6RJseWQJ5lua8hW1rY
I1o184orXDJYOzNywXIIvT47O7Ssdz9DYcOpf+qvnTxdCt4Dt4HppykASvMOHPR2AQseQY+l4YU8
8tq1c/7r3Q1Bf2DuCqWA0DCJIgpMiNDoN5dKmznYOLgItIMF1cJsFA6SH8Qk1ZI9wx6nzG2Em7Uq
HcjI/YzEHRv6wnZQtmu54JaqBeXUpw1ShS+n+Stf0CU0XFtUzQxKI9txcqRCz0PC3i2Inwguh/CH
OHlfszPFePKQCiv5selEDszVy8M9eMOnOYSRHqu3YBSclGCA5KulDrKIYPyq8I1xBafOQLV9mp+q
lS0yUiuwWRzfag4roHHkz7En/6/9UwIJCaeKyV33QqiViG1/0wum8aTlsropUIwxn6yW+Mp0ULKz
WhHHSf80az3apxxq4KcGcbm7T4GPQfKUJ2Pqn7uGv2bWo6BeiEIY6Uvf02GI5HGUQL7e0CXvhXyA
C3twWRVkv8W/G+LPgqLlfcFeUp+HNIAORW1q7TaI4iXGjKhqTdTzCLTzclqgID7JXAwHgLY0kjWt
9tltnJtsXLtdtB+ElOXWljCehdFuI6uN3ip0oLk/c+e9z9tcN36U+kzYf1C/I7iD7henOQUH73cq
WgIvykJWiIIbu+P0i7Sj/NM78Uud44WdAktK7h1CSq43dW2QYFCacDuH610Hes90hD4aUAQuLHH4
FIyC4793Wa4nMjp0kGAhfapsdYiL1E8GMXdpP+tLntlkwAtRxNUUzjpISzvRZIA/gcde7vkik38W
YNCidKlz81LSZgpgGak7KadRzRhoWLrTGOXqV5jAB//vyepX/TXHQVUHEBK8tFfWgY6tJtf9jQ0F
6jVP9+tFlh21vPsiejyuXPNPxJVY+F2lvXMl48QxX3H/hgM6whXCVZKTlOuKQ/iUCrNIXN1zHOAc
z8Lb/2x2oYthPw05xaR0LCawbyNgLmDuFZi1adEB3HT5yExvHViRVFFR414WpeokN7nJOP2pSokg
1qHzlUVtfhvQ4KFEIMJo2i4KnP+zClC2LTlDd78GuMYz5sZBp8sVSUR3L5OumBeQjOYbWPNlw89H
6zVBJWMZAzV+2rqkccUtUd/hTgFGNlNSkzvzbyetf0i9H0++qdAV4mzs4sZTgVw7AT+Rr+Q4KCrI
NyZoOPoxP+/LMZfad3o39QBrl2A+C5TFO9sDn6GHGinvhGOfTFvjPmjeLuSxBgDzJuseXL629qR/
To3Ff7h9GTgJYiH3HgGYi8AuShezhJpe4UqBQ2GP2A2dm5+FYv5jAYOtqGQ77EzOcj9QTbG34FC6
N/hmPkcTVjk4u2BqrAzO0ve5SAwAws8ZMT/8JPb/nc2pJ2DVxRVB8kOoRDUnewk8DOrO3IDL0E9x
VtE+u9opyVpuJp3kt2nIdvDeYtsoOnDmFKHRp8iPTn4juWK+bmTvat2o49Lo6gJdYeABG/1W5rKX
XiSveJ7/OfBGrohOKVFlzv9akqqrrMgpjkTb/1J0QerUI7Y1ju6m+pAaHn7ZZT7hCkvttyFWPSPZ
amTQOWrTJvpFnYqC04/mMxAAXcpXUzg5qoJlHLu4l4E5ckHSfvejr8qfvicULy2u6P6aet6cTzJz
ksV5MMkq5Otzp8pKZL2p+bFmNwoyA+yauywBe0+9EcP9wdR5y/jgKSwaVNzqRmAIRdc2HwWFvejj
mc3oCQN2u6skH2tI26HStkfKzangIke0yaab+4uwTDmWCWK6ANvStBopVo2mX7LJ7kL5/30dOPar
8uV5UDIefhzANiE4+d+K+/VJ6OXokLFY/j4SYpnHaRG92vRAhWS0ceg18KK04IN6JOupm06Ww3ht
CYUNti6YcOegu9USCo/B3Mrhu/cMwvCI7vuRx04hrB+mZ54ZWj3wEJBJTz5MgBstgmzDMr+IKP6B
+j4xzt9gg7tcDeJi2N07Jty6g+1Py8NzuErdPgZ4ewnmzsrbPUOVHFGhDgEALRwJ0zUQ5Gzv5G4p
CCBL2tIeOIrdeESqZpWsbsYS1k6FanJxdaC0ema7JVc/a2tPW5Q21DNzUThbL4TSdNBkH7ub3NZU
8mgFTH4qJ8DFv3QJ37cEoiJ+OKXMJPC/xLd7c+8eKrDRVhc9s5GQm0Nuwf+DTclVVdv1yzR5yxmq
YkQNMPu7Ko/7DKPXiKBq6JP9YzNHrWfSw8omQRdJCQIqV0VdgdGSnmkzU645uWkZb8rc6tdmBXgl
nd4soWCccLpIv0c2j5f0uBuOHqtZ9bx1waz0qmp3qiEd2ZZi9W4l1vqcnWhJFiSqGt8qnZPCZJmE
kBxX6O+0ZFDaa9EO6OfPSGUN7wDpWeHs/NI0hN7J2JiKDjjA680R8yEFGMp0/614GZyBEgMOlEjy
n8EQjgPzUOxiPnHdQi1arSN6KiQ22kqsw0SRBj3FMMIQIdQ5r0eGYU5OVVjXr+qgBXGI3BrI5rKx
Uy61TPXx6DrnzRSXuSnlRDGeCgTnRLzyEm3kTNeiflB4a3mCHMpc4nLTVdcRAlJAkZsZMXjNH5P9
kYXUSv023O/GaF2+w6ArGuwN3q1D9Wf3UKi6cdgyfC423rAS2hiRY/j+y7ZiHgYxyZC2bEoFLGHm
27Uu9bUxeG9kP5skve3cQ4nu8kZOazkiKS8QZLx/QjGFROlveE0HSKCIKdjXBiX4Oo9cxD1XLpkv
LATDtYqc8JB2nUD2hBCzGz9ycWAfc51YBz/0+Mdbz5TMoMN/kWIsS/L2wdCSBjKeRIW02NHwPR5u
NKsy0vGsUhWrD95+PsopCM1mvSwcirDsw3xVEovVamMA2KihJQ75y6yn4x91ShdHyjHqupq1uRyC
hO9Ngx3McZ6t9OIn8lxopjcXlXuG9jwzzgA6Vt1dJijdUWao6yjS3xG5OyeOdyyMhe9u7Jc3WZQ7
PalDUYExYLR3+l6S+rM2a0XcdDftbKcGZzUBmrmVXsN5tDbPXukGgBpF7Z8utyDaPh2XMbtHo6TP
3fLx04NxhH5rvNbk0gsI+S2S0rbc2dGc6Ahn1YrzaoUD23rbgH7UuDArJhM5UXg8k722TDjQM0X7
58bOWXyfx+t677ePi9AhzQU0mZHACzbjtOvAFgeNKJ19ehA06Tt4TkAwfyuUVl7dwq9LGF80YTHC
C+qTakN7ww2o2lyvfPsh8IpXcrBgo/MJvWubFPrYPlqmbkHUPy58Y35ftN8QFFqp5BPX/tb0BWqM
qmG9PcEJCmze8Mn0inhDM0sVRV6UEsTx2bhN3ZFX3+pQGp57QIwW7n7yEw0F0ikVkGegVl4eTqoF
PUhMRfbvdX9y7UJ3ns81JWrJtzI1kwY5Nu97f0MThFHtaVTHYoBnEN3t99MrKagNJTBDk//T083c
6Ykaw0eqekZhmO5i1/C85/1b4HT/g1zkb9NM4iYfuj/mpfN2vyhSS5N1quXFwxy/VrtOQJKoXyvp
Nx41+tqTfUsh2oZpMvd5qeDO8fDcERf9zuiZ5pxAYJJDzZEAdwbAzSG7uK4HbFyxzX/qoyc3ZALn
q+VGZC+HB0o0mWKC9QPkUct9JTQYE+h2EecA15XFdZv5ICz+IO26DqWCTC8bVVzytBeZmDJi4J5I
+1LAuTB+NpdHmD9AgyJ/AqqTG2lsyNLhRkjt8zM5y36oCgmhpwRlbPNPzL2k5rjef2lwfdN+DYml
IG45IJZz1a8FkYIAcXWWUh7pY3QtxY7FdbY6conjJe6mDy31iMSl7imzBRERRFg4l0XxgfeKc3lm
kk5qNDJOjhfMnKp+v6uRDoUw6/EWyNya+piwz56Bb5qK+618op1tbFt0Jgxlxj3Sok4fdAa2Jb3K
sFkEw7NaK/Oo1vDQ2qKvMdaYQkyTHQxEm6P5jM7y72K3Bvm0DqEWmr7sqO42sue7hFAGn81VyF9O
FJU9P4cAt3QSV3cV9lJmnZ22BaN8HpTszX92lzAO/WiD+j4lh60XMlEA/Jg4MyeSsnL3exNi9vk6
RTuXVg9b6reikHhsLrEQ3gCXMeWfpVa3ZLMFttrR9T1Wm1JAQXvGh0wm7mFCCc31buzL299ywJ2D
tl04h6LFMydRrG6pC2Ed5jymdI5GQac/Zj2fKArcCmA968I54xLdp3RSufNGbdHosx33Tt5IdwZ8
TN0mCyin6aGF+9FfsFPxLwWZmHWLMegjQy+rzibBOUia6Dwc1+jgG8cuVGGH4kQ1fSCtKBOHSk1K
JLcm1EGt5775aHPe3peCWu21DtDv0qVCAJI2quO/bYaisIm7vU9iY3cl1ZJJTkN5eYlgRbmfOXH+
ycmQC65KH0zkbw+VjoIG1pO/lhBm6EnkFCx3+tmuPajRCGJMDX5PZ/JnRN0R6bIZMIZ0xRd/uvlh
A78CPkwuHzhllSfzpjAVn4mL9VqeamSVYIxSs/zRVg3Ah826q+Amcx8Bua2ag/0QWnAa8rBpnMU3
ocPY9/7TSlLMxWfCLyD+nYsmTmzHzscyh7h0b20BkwFCsy61RtCKI205U/z1IJ4ijL+g/diVWLXS
GkUPSs1qqZ0WrpGiw1UVMKsP4AiL/q9zlChWnHh+DYMLKrPlmHEI2+lw/oyexHnUVhrF4bLSzCha
uKGmgeTQsbYkNlxNb2MXJsFIVGXSBWTnnpxsRxi9a6kvStOFb1oVPwcsNJI5nijWeLBUCVuWX7k+
3fNF32D12L0GqO03/XTROlZE/xbKy2YfSVYTdnAxi1cCRAsy+JgpOZhA9QFFXlRz+iyAe9VgqkfF
drxSIKSgTbkkZtjA19k4w9dpuBE1B71RWCM4OzkH9Wb//Qzw9kYAI7K34IXxDS73DepZFLKp5guC
c2QGlK+iJBI+051t8eI3ZVfrL1ATzrMdwhpg99USczfSdJRDrvM8zYojiJpKcJ5ZmOFCdoIZaNVZ
xdVdkdXjCe5l7FtBK8yPWpyohXJpqO5JVL3z6U4T8T0vaTiLFzwanIqgEveRopnHCjswo5dd52Dt
cfyWQZgCXbE4dmxtr/r4R7kkDFP2Fx8dH+nJ53bTqER22I4A5F1RNO3zk8hOl76/YKoHvYx9DY4o
B1TXTk3veD2gvQEPWquVHbK49LmxcL04dQHEB7hsSbb6AEVTNLmbGdLzRbu2LbVd8R36eaFMlFc1
K6apJyE+eTFRYtWnXcU+fVkWld2XMk2lzrP2CLWO++BqHfTdWcOmPguHv67CV751B0YvUssnkhDj
g+v/YqAKJYLqf87vqDNb1WRKGkILQMMFBO9o5UzuTPpplIFERFEWC9YsH59zofbArXenJWPmAF/K
JMau9C+6mY6eSoMwk6Yo5rIVV+7fdwvvYYXnHltLFrQNyKrP9+srVNmzmxM+ZOx7W3WGT+Hk8TFn
2jFTUkUUFPQ43HapubRFrAKE3WSF22SquExLQFaw51OMH0ivWd2D4lFFlXtu2Yq87DYb+v5CpRWA
uZ6Hx4XuEVp1k5F2eEo40y5JuxvrrhNQ6QRXnHZAw5Viv5afBoHGTxn6zl1IheRQRF3pbvtMEL7I
Aig1oRcYtfHvXarLXmt2Go0TmCBQ3PxwQO5C4jTgEGQlb/ZcK3soYP+TP0VBJTLlr2G8XfjrJVHT
vA4gGexL7zxAsNPgkg32BYLk0/EAYUskB3K5FVv8fORBlrbk3yQGR2IOGa2PAoFUPoiGXuvX8Nhn
KIor4xAzLR59nO9LAPfVwvyepU2Cvo9hkrf9bPOUr7YTDjocZ3LIChIndAcxq3Q9uajjFnwjRZlF
N7cn+Tn9TkWmAPc5QGx5rxDp6i4KTkTCQ4gl1rdSzosQ27k3pRRuh7IYlZUI/91SI56UZ4TJ16iV
ET6BeYD4Sk2Af/uv0Pxuuh2pDit/xtSc5NHvkiuYnMTPtd0jUqIdFP/ZkAob3XbC32LEofqeUsNv
tKP8D4MkYn4FztGT5/jqadX6MIpyr4LaamJGB/RxgQ/VmZ2pwR4rtap1NdqvgcqAIsWscJaRuz1Q
E94FZxydD+8c2N7IyJktK8o48dlz6f25ocDJIGr7hvFtAYMGk+FYChGX2ZLF8gedc46PgRT1ibqP
FTpOLUbdgWqJqa7Aq6L5ZQdpTRBUQdBAghGfnqvvW+zxkVfxqdggOykq7Ql4iBPlCJAUaVGhuvoK
LgCxDMe7X19OmFZlUlIcMVpnmK26MC1LrnZG12fYcAbBHd1J3vcaxDUrrvze1TstoeDX1wUVVdDq
tfWdJAlIZW0/fTP6feujRvhAOTFOzgYbnz6aXKoc4NFqW0f8820aNoAfpJ68nmh6RSySvlfHsvlY
amyt+Z7hFOF2/6N+fCSHyQLjjdO0PUR8fj7bmPqxWUWKrMxfXVfCDYcITfmwyp77+boR09Opuvcg
v8RVpnvjiTFROuyHxbIUY6IFLumtpZiqSEES8l/t9OB5G7hbnX3zxUScJ6paDie/Q2YqfL1rda8j
5IRdMvAoh17tMkyrOeNsSN9b3DaeVu2xoezbzG9q7AI7o/cZJXWRj8ZAWkWv9H6p6UeaXVU69IdO
oKWWbrKM3ew+9sMJWfXqwB0O7SHt4eL/Bqn8oGgLMHZ2mGN7wlOw+gWFL53RxLohlPkwllMuU4ya
txf9rLWNy4OGbDwbE3sWHgMsrYX3gjcJDoQQdXnGmblMUWeH3m8GrH3d6pPDX2VElldPX92IkUL8
RhODMCUVoSivXMLduYbfmsUrAbf0A4Fp4EFxrxxnS+uZqegydJUq7QEdu6JkrXMeWrIxqmb+IOdT
gAtPZhr8I9yj+g3zq6qx6oIdQUY+2ZiM5YxO/Or8OEc/5Tg4Et1llKkWxLIr3b8RWxh0p3KwgaU8
+uFYL/N8KsrPN8EERFRhmk1ZGvf2Vfb9UviWDGJxmWf7HcjdBE3cw8R8G4n1GTNlsaug10PMQOg/
UIH6/T/U8gwHyD4CCM9qFyIBHbT5t3DGph6hBkhBGaQoY0QelC/nqwW76WQYlyzPJdi4N5PtUHKH
FWvSb6nnCsJBwApdM3mRwSAAy5r9I67KS9ppvmT9uWHrAWGvuoM7WOyklXGCFonCY5C8TQeTOk8+
k5EMEkmV2RZLT+92nD8RAFY9pyL8Pv6d6yfOdnAtxLm7OcEaYqr+c8MlqfprKQu25a8y0Ah86WEG
xkRSiH3LpRaOIhvh4XztGNTa7/DVCuBQsbH+c4tU99Shr2Or+A4Uv6dWeOuFlXQ49fns1bvAnRgd
GLPfjcJVnowr5FYdNCg66FeZbPwx32CwGhLbpLbYnBC4a4gU/H+y5+Ey6QkmNomIZMFfvotE44ZS
zVgxd7uaKSAxR50Myv6S7ty/3SN1cWZPJ5iATy/PXUCQZOleSU4Kkja3hJa88vBuo8APFPxNPMj/
zA6OpwbVHPda4HiVnNJMGZoMTO3NzTb13FCMQ8IbT7Xv1bvvVnKXL4VG7KQqEIgLL6PgApx2TPXX
/VUxM3qMNA0WZ8us4ZDkJ5lGBmScxDEWUNXxma5BkFBPTjrZg2xOMAcjxD10Bejcv5KPxYOl6+mu
FqCbC/G/ZiDWx/QwtM5neJpWSsSAXg5aZyws7D/zC/ZEDY5KgPb+87zOQ7iXjSA/jSPkODHAbVI7
qdzgb61d2YsGAyiq+jA1zfNczJUcgqLlggshV8o6axXiAdAsrONXjd3FXzhO4ceSthphaqfXD2Nb
L9+2NUJ0D/cmP7Pp+riRKV+F23OzDHcf1TtvKejPrOaNwEQz/m39h5zF/7ACbLyDK6U7le7SVa29
kp9aT8UYtm1fgL3GTjQ5OHAF2toJYtl41WhLoz9xR2dxuTLBvRHgWU9SJSMhmRykv3EuenA8JNOu
Byd/aPJH1x+rZma4bkJ6rDHfbm0G19lmSUEr2psIkPSBHdxGLAYT0xTmDEywhME0nHxmVTZapYpE
sVpT1Xj6T3nG/C8MXI9iCsmn9QDssvtxkmftXHAyiYF/FMVOaiybhcezMD0hpiQtamlmeHj/72ek
0PuVkPo2pkCVgIznUiyWXpjbF+G8bm+4uocuADhHkfxyxmvIGJs07oH7I7RsFBzBTmcylsqC3JFo
hyTBubqEB8lAHQhdjB2pFihWUswtl83Bl3QDiyYi1PYCpXGYdoVXL+dNZ57Lu1MgyrpZefnkwgTj
Rlo1F8NqwQC6itui667d4qR9jH7QqYfWwSyo8GvhrGQayK4oetxpBUPVCelbXK8urejxJasyPLDN
tPekswhaHAOWHNIVPgUqiqVAecTN85OAh6OwK6T5Qw5Y5rtMlFtWBU7wCF8c/pY54fsUMlvcRXM7
bvrTNqf3HL5Zq07QOg9+tglKAXNVW4ggxpVxdiSxXZc+gHbKmhe6OzLZHQNFGXUBiimGhdQOCKTi
3jyiJLPnzCj3OiHxXoC5TD6FLx85KgM2Lioaux4ATCtqudwNGMBsUVMpHDfnI/+PzUVNWdwkERVQ
qThUTP7SKT9WpUzX7uV88skNKlUUYD0PKXzdz+cqJ5Z5SuHzv7I2Wea2DiIiRqY3iwFpg8FIeY11
u/ZNrenvjFtQlAAyJATLzMLsdk0QWVl7vCh/mc1w2voTERcx95MXcV5nzrsUmvsHuyhrdXBRroe+
zPLrnsMlqzV/YJovaGn6RqtB5pzsoYFO3sYHFks/RllroXdk79KWD1ot5tEh8rUxgmw7UrzGPQuv
NtZ2hXOu0kVkc+sBsCzDAEy4LBfGmKMbaxZIsXeeWf3ab/mBcPxu0PZuJJUM1whmsxoSzoRcnmDY
Fs0Xc3NVYkfHglD2SG5SiyAYHz+NF9/BitjId9+CSIKcTacRV/roszRYYbDgcUzVOYzW0gTW6B7e
E54seO7F7VehvSdeutuLCwhEZeXjvonWPq5mT00TAdMbvR5l19Ykv7qkLPEeJKPbMMi0McKhKDLX
0Ouj5esMRtKJKrtXpTJNSCug66c3L06GNGFG/Dc+Fr7HBGIX1PSelcpIH9QCh0KzToWEQ8ti9Pvd
stDpki12F1E9hSri0Qs+89Qjnubcp6sjEMSDtpga0Jb5+xVCPm1d5KtBF+GH9D4EEMI/fwVg4fm2
+RofY9CRSnqRMAH7ZOZvVNqdG1+9XWiZiKO62RgZ3HjnUyWmmPu0BwjfYm0LgH6KTw2RpbXOX7zl
E8ZictTJ7uMV1ICW/NMTj4koTb0slB3lq38wmcHlCW6kz9syp9zob1oMV0nX9I8mM/vdJ+EtP/Q=
`pragma protect end_protected
