`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
d5Zmj3hyPAcqEti6p86H3pl0HJMug65sJ/2DufB1p8qzicY4BXX8ZjWGRElVsfOKzsr2KCY8N2fb
os+FynCdbA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qQ7AVQqz9NDNpNBdXK9bdW8nxNO5fZiuJ8SoJjshbvYEO+yDAJ9nmgMTQws5lZWTfIfWacH9RZB6
NaXR2yP0fWvl9M/UjjwfohyoAyOd5wQcxJnhXjuIMCWuhJIpoBhM9xLw9+JJ0pyvosCVHIeasE+2
5TXopJrMtch1O+DUAUw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJn+ku2zzfUeTU3rIyKyBdyofDpzo1w1rv6pdx50I7/w2xcio7L/i23jb8hO9Oj9IGazlSCWi1hA
iGUnnPF1BvjvD632NmU2kzdfwnAsb7z0jMtI41Ynntik/8IpCV0YIe7eSt0Pc6O1i3lCo/xJFYp0
DKPZmcIOcc0OdfAbmpD/eD+w2N2TDx1YTY7qNWDwnsNhtgs+QZIgjnLmhrKniePFSJXm42EKKJc3
1wl3/GpbEfltSQ5YzWuQTGqFgH69i8fG/pUzDm/tTtH4lPlXRfjaI5KxxpZa1cfahx5mBxslCL9k
aJL4FxBpz7nFx5tKeEegfB4D1ffIav5oT7Z29Q==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
tri2c3H0iHtN5V/yK0O0lDzKmG7e2HTNZmBZID/3cDYY5sxqJeVvuoorB6a6ihDkbhrWlUyQQdnN
tLmNYiauq3YAn9kTX1up8QovJQ+ZLn5ynW9nrC683zhlNV8iCMk2lnTAn4IZEdOasIH++wKrg4f8
ouT3HRFAt1dD/RVXY7M/51t2uog35xn7pMJ/etpulgmT26PDdXwMeqpO+EAQT1DE7fY/fm/4HtP8
Lh5KImFrrQ79d2yK/QQvGpVFAHAGh/jXq2FJqEUkgyNXo6qjMZJz+vN9zaL/nsfXv9m2uZSW1lFL
CvW1JmKZFdIWjTwrCgaLvoF5OxbJ4vFd1oHhRw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Dw3NStz4urCgx5H6O34t5gh0C9H8xkUKp/LY2dcjrUDocGPj6rFSgpdvvYD4yRVdUAv1w16+qnlh
Mza8XJPZ7S+A9sQJzA02335YGZsvoq2WrK2TIAKWMdyOYC3UdiPATr1m8Nx37Puqb3/vHPSaZV/u
lX8CvizBV2pFSDMF8efPgKG24eU0LbEmRaNCZUBsjH7hhrXh165PVIxRQ0HDE1mWbVv/kWGWjCju
D68C2vbHAYuemZwogAIfnvTX6216pm/QdtzgeiEgAwiya+U/uElGyYEDG7kALz0+E6kuEWaENOiY
3JblEPtZ/DBKew50F08qLdI14sA/OYlCOOiduA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SUxYKzbxlWiQXCkP45YxrZihOzRzPjb1t3il0Nxa0FINEDnXIzQ8q26Et8wxpvYyRoHW54qH4IXY
YggumJfU94iNHpRaNpUbhB5y/O7fHL+j/HCeqGntNjq8DO/4O7rSXg7cpNlw0bMa5SJefKqHIF4A
RG1io5tEvTk3Bob6Cds=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FSsk8VGUDHy552BAcCQpYKeUZACCw1lvfwnuDYYGJctMsn6t4peO9nlbm07WR70IULjdIvLq3w4q
MFcduFDcn7Wn6RoZ08UXzXS+q8MJkJlcutjgcQAJSiUm9ZyeNmSe5tR/OUU95wZqMgaCyESUy896
LUMrCuEDP0xlTleigM9aUtz1Xw9Bzl2gO4kcDFOt/0Xa95z49To0//ryfhUYUGDkptprJRbUfcEY
T/xg5w/HWe6Km8jmnAyxi9wzT3NCJu4esIN1gzwFUaZ8XF3cnHw4QzsROFq9UOHmCjs8hiuV0Txm
mAYF2krDEmTvkp0frLWpgIYf8Rv1yL5W47CflA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
Tji8aM5bCfQrkdfcy+DKS/FP1Ez///MeBrftwPE45uAX71Gwzz5J7JNGC1j9xQpaW/XEIO2ujxpj
gJwcJq9VEjTVFCdN4GaT2Q6K4Hqj/cK4unO8N1lkY9zQf+80GpL9uD7E/RHc9VOkQDZYUxDCgSiv
sIjysbUdfnmIzMp+eqkPopDb9j1Je0lEgRtq2Wytm7rHwRNqoLEOgoQyDr+91IipYhFwlBepAw1N
VWHnfYaUC/BkjY05VtebZaiGVbfMifu9MYuBWMpdd3wa719jjHdptqlj6/qcCUYgCrOhsr3c1H+E
TvViOOXiLTc0qf0fturXoZFmHz4ZFmeY7MhSu5dK2z9g3pJUc5LbSefAyAJtKwXYweXgnou1bOoy
6QY8zKk0OYciXSWOtWYDpvKWMJK/G1nKjR3tIggehW78+JylsN1TYZ9ephAOAc1gEPQdKPblYQCB
fEaGPpf1jYhmDKssBXqarhH4FmMXhWmlCXlVRUfQwQcYhuQebRYvIMexhdxDURj/SSZOV9QLeoPT
VJf+3LyLbUt4o/quz93l4r/zI1bYHmluvBXPaTyhBL0jDRfXECyR81DBlUbmW8PFnYoSSbmZ6Km6
D76E3SOoJ9kAJE7pP4iwf6GCyhbIe7QxGJs6pPPOHI9FH38jM/fPPkBujuaVHsM2AeZBJbxEExI6
2eoijq/IZVkzbdTXPL8g3gGsvBQNkCpbimvJcb2Ci9+n8FY8nKbW7SPbu9Bf3C9yEzwoC3+xy0zp
BPPj+2tINTrtmSTDnq5+1tpqv9WDg1WAL1YoePaeXNrWSGR9jaZiAWP3bcAnNgo5GWSVt89GZaf0
TChNW5BL6P1Xs2B9F0LqYNNNN4UqXwBppmi2GN6vVzib62uK1bESXsh0Vc61yPJ0gy1g1ad7E+jp
vEaayfWgSPvOm76L1GhsVuVJzhAEkeIjMH4mJ7PsjizOC37MI4L0UHW+v/9G+F9edqvf1y6G/Isc
RBcB+kcBAWb90ReTA85xZtbzTQYchrNM59YzNyP6B4J5CZJeOj6ebVzPoh+UiCxGPgZv4yaMukKs
z4NzZigB0EVu557iu/WQwnwi031GEX9eCd5KVUoC1rsWH7EmlbMgeN48pQV1nMEFqD5ktfN/NwFO
muQM8ozTmSbW2KjOwsANylDp/VCkIkFG+tzBoq086QUo1hGfghgX4CvDZScjXw0VLSRGu9F4HN7p
MT/VO0BAYUQTiZI7UwNmjyJE1zUUKGah/S6rvYuCWfi/v0ITsu2+naHYdSWNVbmOQmzOHCyALVw+
XoG3GhfBEWhGySxDKItj/c2sfOq/1phGGz2rnC3IRXMD1DPHHX5I/BzeHlFOv9+QvtGmWm6ep78F
qagHvfpvB4xqQ+AjT6srflbhHwfN4NsLgnlIzJCtyciI8VoVYo+mez4qdMD/UBA2Nmm/qUY1HO5K
PvU8V+Sovn0T1Gd3ScCUCMg69IkS5n63PGoXwJjK9HlOJNEE7zR/gK8vTWhnMRvy7nOAXH5v52Xs
+AVsGjYW5eweYuYJJ1yOLI4GTTXmPdAZUSz4JA4CBjbS82LxVUlhsbi3iM1NoM+5lyPL1kDypdiu
MNUjm3wmkUwVfZXMqiUiPT2+uu6hXKteVyByTbdetcLzVjiPQ+gN1VBf/iOdR8uicSBezTVT7tgr
fgZGLZ6owPmmoWXEzx/WNZQ7iDgBwFMbtXUQHduCX61cG7NAmKiHY9cN4X6TZ/R3G/ZnU4nf2jOh
OlW8pC5LO8cWl8kKVsVJmC6vBf/PdRANorgaEMmgRffAgD5RkeGU+UDkqeivls8HmpUTDN1o+kxJ
JxQaGdr1l6xnJ+HN3Vlf3Qr+Iw5NCCsccnu9JstdOErbpylaZ97p9T8YwUc9LNb+r4nzn9zbgNG3
goo+DvYa9Rdt2XTAOHNOJrMLFPgzhAxUNzrbNm3eQ5ohRI9jRxGKrFPOrqFDsjFCYVKGBDVyXmG/
Gj2qH2qabGbmt/RF7as50nDzcjpNq/EN18klK7N7q0JINpoMfk8YLtpZ+QsEvk3U1oxy7rRXKjj1
u3YIrfd5jq1HTdbp47iBNquvnJnKFlMrNPvysT+/9ynvJFQyLdtT8oyjjJakY+LvVxPHkUd4ayO9
ozHiJtSjJTgEY6/zOz4CocppJ87L5E5dm6qv1t8NSJtDZ8Wi16NondbctezsWEHfq+lmVqPo3VwN
VkbmnUgqHIUninO16r3+isbNDVTNvkgtpbPLW/QyBtkNSoMvlLfiDbC7rBbdcMadhXWTTTwtiv4J
Bo3DpRaHTvRZVbBqoM3wW00led/UL2Xs3aXRNQewasAYB8eQXA1HqOWqGYndvLlCh9kazCbmalSD
HQAZMJFay9IUcNcXqErRrEmDy5s3n9Ct5j5qchEvn1PjtrHGhj9l2LqdXCZSTcFDh5KpJamCNrPe
FmCYpAyBVlbG+WUQV+siz9jnGjvKCIi2QFdgy4x7CjoQ/fWqGFGWrh57qAXqF6adYFKrSSrsbLG3
7+3VvjwuVGMV21wviuccyQ4LQTgU7loi1790D2+GGMQcSB+dZLKxq3D32Dp4fFwm3OIklI+hatPI
qinPhJ6ei4x53890jZwM56G04qOiAkzScpPbiq100w19shk4nYsei9lt7yKO9JHjM1AcsALa3XYl
b/hd30I5xI1rp9s4NDNetwOUBqhqmd5DTJ9rBjII6nrYMearjt7cp+6XFnqFXQGZrL8JlEZ9SmqH
FCZ6t/YmXWV+AjTg0aOqL1h8MH4cEjOu52BrIoNJaDfNIcduZWY4VL7JegDUaBiQbhaUwHB5l13W
gPhapIMQlHOD4/jvLD0LRzAicEBlNkYCsWxMzo4F44/43OTCjMiikU4k0gIxDxdweJ50ofQ2uMDW
gbdVQzF0U68DaUykgK1B1eDl/UG71n36iN6EPdjAu2NlRfrHh8j8L9sQ1nwG7WahGbAqejRvOqLU
rn9znO45/uF8mCKKcAYdnhrlv+IQq+DI3+BD3g4kkOUwgqL5BHBFhmT1E4Qclc1J4Qq9CpkfLD8J
nv7AVA/sRDedp7QIihF0iKzgKZrQ95vni6klbf6/IcoQeNS7fMXXVVt0DnieEdr/jZL7o+wG2ls/
c7QDiKJ06ccgZdxRgBIXB/P826guauksLIlZRf6VnepYAfvxV7iBnnfzyfm4wlqJ8IhNsOc4H2Oo
gz2h3ErEPMAla7jeeiDIT3S8TOpTF0iFv0skyZej6v4pcerG7G4zQYCdA3l9qF3P+pN4dmXDcrzO
MBDug6Ek6X45rXR1t9vV1nBjjWyhRilkuVXAzwH7fv2TPHtmB5TwLM/fflhX0n/sW9ml5uNsJsNd
e+1BlCLhWxfH5NCVv22iMHDN9vnRY+WFdW+BtI+KPI6GLyMnE4TFZuX9zygIRsZTlAjsrSp0loBd
2aaVYQ30vflhg9yRcBMz7oJketpZPQ9B0Du++rr9A0H9/Ra2Qrrvkl2f6gDKpLSKnYWx0XTjm6c+
QnofqzAfn8W7wWjvIhZW7WEW9LnOzlXPP2aBZIcJqVKPPLOAAujRT2tun73Zw596AupCwNwDDcLp
5FbbKqrdp2Qs+sKIcjFa1jVLp8siEgygrhG/QFG0WoJ9gCPo2Kvc9yRkAHT+BuPf1SrOGRrVkVpz
TeWwsgRK3s7etEJD5Q0QrJYAvWK/ULWlMrdTe0Nwg/yod9bjY0F4L/eXYTM6JNBYc05JMmGiLNAh
5tr3X/+My/wj3SFMdpyf3fcu+Q+bDwww9wFRCyNsvCwFbkuw0yMmnXTBJvsjN0N9+WjnOLsl7cAn
jEKzYR3bxhiw2MCn2iL1WfMudZqKhaQTPTjGoEh1iiN22O7UGyZO+yJMkyY7hJy/hn11UJ/sZklU
zBGvJuvjPPzEq621r1y+EQIcV+QP1GBttO74Jtm4PEW/hnzlIwLhvQdachCZodPEj33XSR82y4W4
/udafUP0M1N9xOgImSL+YfsHN8PWd3OjQh1gcj7jNvB/VqLCJXEVspJgykAg2osUYjm/sA5FxGBa
bdMTzbRhCKD9MuPqA62o1Ajfh/l3durq5PVxbTRZ9jqg6qRCHGQP4wgMHlgiGj7LLnUIT5Ch1BaS
gPkW0ulvjOwZiVbsCbDU7/ZrDrFQh05uQo8/8EVnIKlCvZXm+Vl7+3GB4CQNFAjtmenB4iLc+nCy
9HVOQlTM8RRUMA+js70ERaCo/Si+u6WtQ+QCx+uBKW3ZmNfInAHxxtWZrL36IAa525ObiVa8LkyF
45mCtbgofbonmmJnZe+Zh+Bw1v5RCoSgaYjp7IgdOKBnrFq3VcbaYM7j940DUrhmjMTEvypKtf2X
WxYp2zVypbZTM4JpTOi19HIkH7NMc4SIESzR7CCJoClMedwPUQPh2JBJ3QJ2zCns9saBaTzJu8IO
ACKJg0PYb0BpbDvnIph26maP4wL5ysGb1vr10vnQ3uW6+ms3UvMIM57MZpdT/BIMu9yQ/lXofLDc
qzIsRku6ySrtZkiYgIdz7Vudh8OhYReU+RdFoH+squ1SFTZTHVCvWO4NQ0l+hX1m8HyAeKU0vH9x
HSatB4bGQ47V13IZ4H+k3aUivEkqSj6Mh24xW2aQRf4ypXwy5Y0AzdGcY3OZQL9ftwQykwBn6wgF
j2nE/J+xSHDIVsEFzMdoXf9GCTyfMW94LAuiU+xOrZ7+7y8jCZc1tFRLI3k7a4FqTWEKGyzY8cDs
eYgiE2HKBlQkwyuYhXH4fTzn3CTS+qx3g+aLpND7pYzFvubRGh30zoxZGRjqKpDKEV0l8L1hiRiH
B6x0Y/s2JFXQqqNbjhR5FO8vf1VdUEO3V57jwqd9Q2shfa3MRVOURj+o61k4eR1NaZ/rqxP4myji
w85cxTN+ItFa/EDCg8LBHShwvzh8XjQBD+bBYWieZNguA0lRaPqCtbQhJZXZV4n2TYmbolXsfvbt
/ZHXS7dqPrXmiI2v+BzPVAz/QmFBziCYusK27fEfEf+KXV/+Ep2EItb6gxmrRVQ7D1S1OrEHqCO8
UYXp9FeQuVcyrGfxwc4o+T+KhIZRZCHmfpccxI+aeHr2vxfe8SZALKdhozdA1HEUeZjbyLkO+Ywa
fzEerHWHJ0v9b7fQJRXfz1x/i2qOfOtIGseCowcxAMI8sYyf7cTHQ+kUzKvD1HLR7+07Sq8Uwwwh
FJfoCdaYYGzvZ1p/FwajKE011VG5Na9tjo9Xjttp992g/rPJ7+ueen+0X3PxcMrjiXWsqNaewcoT
VMNqtcqGYnh+yS0BpEVHa2lw0Q5/6sUcMzZyGbniAqrPoA/bYs2gtNj3KsyuIXa3NRKqNOEV4oFQ
UtbwfSFGg+osVh5gQw+QKZMdjJ7jLp36VeylITwHTnTn6R7p0YKBdT4eyVClYxpKni8YKYGmK+bV
X8rtLJD+R7bd6y+rZ8wIHz7dDYN9tAqtlxydBLqsrWGt3VCy7M9QyjHNs7JQ9H0iFrfpVAOYIgIV
/e7xUfQotQZCbam3Y6tXXARQYzyh9HfVjOQ2ujqtSI0RbHp+3qy2Dd2opn0I1HYBjKbMBdqTur7g
FBU+yngqnfqxB6NE4/AuxwFBYc0VNcWIYKUIb4F9yKVmGCRtP5Om9MUNW1hadYd1Dih/0b8j1KsC
acwSLIbznHJYoSo4L4DDkz1Ctv2JE9/UFq6gO0Lu5NLoq2MquK8C8O5GSOMdSR+pN3tC8MK/J8F8
x4FhszJADVfe1aJAfLPLRtyk6WiuJbwSiWT14/FIWB6CMfxzp3uvJj68ojDLbwR1E1kZFoyZEstV
2iTeeZbVmxZgPNOfREipIYk4vZ467NKWDJFMXoMgupVBKwkmvRFu5Rnxai1X6H8I3kdjC7yZ5JLF
vjX7V6Lr4gt6OCUXT/LIZ6R+BJEP7aAj/qEckNwFbKZ8WZrerWQ7qHCeGOfn2ZFj6PbYM3MK29zi
09xg+JCLULnxaxCyAKJ8EGDYYkrRFWuOZshgi79X1FKXeXppAH7pn+0I3+OTc4D/vSEswsQ3jw+4
eoeAcYOln90exaql94tNpJwodM14ojtzAXlQ8XXugSsafDmh/37iwzklggpE0s8M9n2+/auVqL+/
35Owlc04Aq6pwP7rhkImgPWuuknGmqItb8DK6Jirg7bj0BWpGCNkniK9Vq7vx1jrnincDG2klxDY
jFgGhj+LhESf/n+56DF79eTWmIDrJqKJOJkurXJEj+LxYDuLtsYcsuNeINzuDT7Lb0wfDCH1H2SD
86snv7r9jRdqBqKhFNqJsYwNUwsyUNlkpOEw2F5+8yfQGFIpGRmr+c7ysib8bKBjn0etEgIgDqPy
rsQ4ZAFrKefcUhZKlaST64/+qN+QwF5pQdD/2uisxYW3SjO0DjPT0T4gSFCCzDVbXJSccrAiWf9u
nxHmp+jF8IOdOjR8hbr9omPuN6ERkU/UKYJFQwA1naWTT+ErXgPhjIHyx7mwPsqsE8+Lt64T8lDh
L0W956kKa5eKgr4QyetZzvX8x4TjZxis7NVfcU/ObKm9u8N/0HdxnRjkht8wcQcrnp6piY17iOr5
ug115QNAzPtOXF7ALbubkd8zjxWe/KcqHBOClM9kn2S3n8C7rwTNyGgzcS0x5ndTR+o+APMd2DjJ
0WNE9/StXp/jnxYZXCF74X9eMgTKC1b1CgzGa9XAFEvI23q9XlZ8s00zXDS8gmZS3nCzDS5DJBoD
u94x/hpf9wxhBOjpBUlzN4POV7ApymCRmjcEK1+k2AXM+d2De8FO3oTuyGmtebB3tQ1i6vhoLb3/
M59oJ9ntqHhsEUpT98H0N+XVDhqlOmmXWZ+j79Rf6qsQZc0PMO9QJSkfT8LQQqh5Es1mWS29oR6x
IEjOLIJWbvzvIOf2WwBx9ecdLRtalOxuPekHGmgDdfjpzwUQ00XLdLWiFQ81VT0fjwoTKuAWfBh6
sEHcUmE2UTdgIK4qMxLMbyAFp/F3uNdmESVZLpzaSzCe5P+79XKUuz6tG8jxWkVnIivAhp4MjBZA
q7VMoLTHShNv0gVCokQ5OXR+06wplpkDfJLBTCZ8rWalqeYhSQjINs0eUGwgvvugz2kjv0pKA7pR
zPlY9gms9jAWLTNBj/Nj56EyiovvmiemgtA+8TEizvAWWet0ble8lwzqfkqR3s6JjMaGYro2L6f0
cUCpyVIsllU41YqQ7vIN1pelRIUiD2i9Xvpp+EfaCdveLHf5behKnooqpHbCImi2IMn5QoS6SzEN
1cTRQ0GWf813ujVOUAzFZHhZGpAOj85NaLCA4qUeQGda83KfT1hJqGzg6DHBhDySN3T4fejWp49W
zRxtFFVrhKP1Dbkvp0gBYdZ+3/zro+y+ZxmwcHe9ICMYmtKjoFc1UxXpcgQIGjRKD0HTFZ4KZmZv
PXSGYR9VGoLI2UUCWteN1ELGjBqWKWGtnlYb5O477MRLEWKK5PuAE2Xu9pys+5pe4VlwubttkP7k
amyPD6zyia2k6GTgVB3z94BzsmsJ0WIdqG+BHpdB6HDzML97+BJN8pjBcQJN/pk0kOwm3z9228TL
eY0SCJk5XRBe/dOH0GsfNmnDInY2oU15GCRzGSWN4ySfhY+P7IwYHkmekXYvibYXoK6nQe0+zCns
Du6lMt6ldVCXp9uAzJt+eNjZNAD8jJe0qxaQ6/WzV+e+98o7FOrr/vy4HgCXRbpyasaT6+mKQ2HA
h6Sqz7dfhTZ8ISCSKJm2jRVvl+ECZulZdR6UHZDfAxeZZMYbZniHxBbfJNL0Swvwg6x//Exh1O+y
iILHtyhRF6yp7uOjsJuNXLMQ22I1M/x7FEOnW1RxWRrH5J23zJ9WpTHlTFU/gWNJS6EWtuihFrX1
Fidwp6k+4wMNlT1LhG+tFHqINKBxsagCFkwxbHISR+NkA3uV1AZUvmW6bJyNtnetXLIvu33SkGLR
7icaM+SJEZRg7o11fQii+9bJGIaW0qxhsWWYx+JNwj8SoB8Ze3XdRDEIqVAauh9tQCDunIoPHQOI
lgxoHEehtT6LQEN3GhRKi9px+NBRUyo4f3Q4txWJ82y7Ks3FTU0wqMqkv7HynBrZH0ME9I1ed6+3
BnJZVGXGWvMPaE1r3/BQSiQ4Gg2Hc8Ib0YTZiSSJ5mytAPWKGsEJIpcmg9ZyxAlLwh5TaTeHypoA
DB5eZy/Bk7eVLct/3OohMKHWHXISmi2lL6cCV07PwIVUmlDD3OHnNxzhQnFMshIIIW8XWGldaJmb
iEYSZJqAZTjz1t443+18MvQPf79/OQGkcnPHzFmFV2kPO0CjdR5PYRQLoehOrFZWZXEtpd8noVKm
8k9GtB60nm3oXeaE/QsWXnLR+05nGwFq3L52eV3IAgNulrnW0KWhEcGb4Vec7aAh7n+KjEP9Jn5M
1TSd/WBjk5rDvFEULYCJaY9p4587S5LgfUlAJ0wHE4aQzPL+3PR2N4O5aHtxxOQL1qidahgJz9sz
YfYRVshpZ5Mu7opqV2MivsqUZeT8sNEBtctRCUk3VzZEXw8r6ivFLGzFH20IJpyhsoqNyKTkoFft
XueSo5mWqxHHcrysoaoXnqFWdh+SSEt/SxjYgmmVO8qljYrMzSZ2wn+SI1+0GfN1vvBvW7gExGDg
aRFyTpjKdkyAQtPR8+30HK9Ekc6JOkvRJQtdZwXrXyctlgzISbnrYXYi5RBGqReRORzVVauKmZzW
/pyQqM76SsLe4OOaubIyw6LJ2moox1SnCIDgyOi2y0V9La/8yJNreUmqalCbFOPgvVHAoTG8cy1+
cnIvB8MfcAh3Fhqad4Hv7/sQiCNCZMngBa2xBbdpXVGonw2zq2nzL9lLM5uIzaTiFzuut9ewNzSH
9yagNy3XisDDaprhubAKBR4Eb8BN4OUsG7dzK/oou48k3zFwWDVGkmiBFx09JvZSPtiQk6Ws5LlR
z76N5Wn0FIi1EoZHVHiMqt4JlxYS+7GN22/JgvqEtzIuy+EMR8XjLGQdXulXRKQ0WHq8dnETNqWF
aE4iOucbn+SkFciOV/XekwQ5eV+AGwaHY6OyTCxephVBOp4V25Bc7k97NxcYkADfD0vMSq2xTSHy
2+KAyRqgBhATBKPg4Bt/MgnoY3g5cKSzWKYkWdSDajTQnBF/xK8FJBfNH6ToK4yArhDH4yK3QkBU
ZypJcTfMhMdAqAHecOdfLv+gc4RJycBcg7pUC/KZ64ZwElZgkTUxeUGeH+Dv3c+L2gHTEaLjjw8B
tmZP7nvDO6lQciteMxHvFqzbx1emNEQdTMLWcEqUBh32jdC9iy/eY8xV74+ZtNGlRMNmMJlZuLn2
z1LTzeZHP8MhV2oNP2AlQlVMyrOAGAvJJrEJ10HWo4hxbZXUMVkRFWMnRJgdAAWGidsaT6AO4ogg
+3bm77jlaX2vQn2vKD2AdXd8cYbEFPwDXjGc2hfekGIPXl3HkQlDM0NvcqcxVMuA+n8FDCO4BcJ3
xzBav4vcXhW3OVC2EsRFLhrUT9W0IyhW4D/hHqQ9gQ/h5WdReI2cGhiW4eBPayJuG9TQA/Dm7n4y
6ibz1md/V6TUkXa6JinR5Dat5NUntlfPiYSB4fi8+6i3S4TAJ7Raoj+EW6Tz0o66xzN9fEaOyCD1
CNvcOoVUJ79IKzO0qqEwW4+OWshZtnuXPWhsG5OL64KeUs1kv8EpMUuQi9VV1Cvn95fWTTsQRuSO
pFt9s7L6pFKHyMNfLmdaa3IlIBPf7NKjKQxdhz3848CKI46WTTQjt5WzDxnXH/tB8GB70JsmoQCC
GkGgRnWRZKyrXHPuUCNvNzwJ90rorHe1v5oSHGXg6QIN6NN1cnXx1vNmCMrdEyg0JQT0kmjKYD2H
1mkC3KOOKLiGBFNR899RFsw0VGd6iExFYlktQ4k0ofyrEsyhnwa9+imACZD90YeiS+1WA34d6/KI
tOsmlfuXXr8C53zWxtQLdwhUgZlSp25nma5rlpwayrgX1L5iK3CBC1MTF1lvzmxCHSmxRi/bLPPP
MLGjsjfy3JzOKlTMwud3ACWfPVVPln/Bnt1BaKIIItqxQs2MDFYQb+TsbjrCuhMoGJmaQYdIYIDu
8he65qIuczdEubWx+9vJNE4fxozyqOgi/mPmMyuVUdv8mUM64IbJ2A2t/D2kg9doZ3LISvMaFrl5
r7uUgAkoYNqar0keIzVpvxI6cF7IYqqaRHAL3HRn+mAhtKuKRYsZfIk6J3CLGYK0uRsEchm4fTBS
LsrDQaX1RSQfEYi5P1W3IF3VRKQzvoEqK69kD9VOBUFA2wZ9Sg3qzUhSZrUFUtBBchtcNI/Zk+iw
9QdTCp7IHwvD3n7GTPC/GU4m9sEhgWtlxANrSKNOBSjbrvN4TTKw+tXL/fXnOiLu6IwqGYTIPlzn
YMuzvZmUkFeqU5qd9rhSpkeVF3N2mOvLdxfQMaO/52DY6SVB81OiFk7KXCq0t2KgO1w9V7L2tftt
lxHKBwHVfXPqVi6QoRPn3Ys1iHzfs5WYrobacaU3Xx1lQkP9DKR2pgCTcJORB81jCNEtDGGgnsWX
SWKNNAJXkb+Td0ZsKcnWgekO/0mLU7P4vicPnaOKyp2cCq90brldqXdrDIWpT8WO/l6JFlseuQ1J
2EdfftwN4jH0ma+5K7s2xouGgNapQ6aBmH8w9SkaTPi1Msju1AwygiPuYCSe3ZhTyR5n8MGh0BNj
TFJOodI8wjiUHOJRkXH1MevYdgKfImESOstSvWwPCv8AvPzluFM0JaqV/2x9p4cNhct+oxVrbEMB
BxxyY9CPXPx8X5zWVE3ykMa8LJETf0LEtWIcoZCpGyk3nC/6oTMokHI3c4JHqFr5tC2eNlebPOfO
H3BBucoGEfxWqCgj51mn79Fxv0koP93EAM+RJ9Ln8EFXK8Ag2/XlThTtmiBV5m1lWIQ3CLAZ/Ptb
BbHWg9o+B0O4t3FgH2JhhEgP26rn9tk+LLJJved6NNmAopv7ru3xhYRvJ/fTIta/MP919Mp7fLAq
JM8Kr0k/FxdupbIS0yuMKGuXVrbgltqGjXJOx+2mZlvUm0hn0az5pgCJB6palrxkS66n6Yia/o+e
PlhjtxfFP7d3gJl4F0PU9D6d+joAmANJ9c0YhOLNGKXY72LYPvYoB9oCSmi656Ne9d4/ehChlbU4
+S4cIT+9j1Se/apkKSumK61Lcjif+CWx0ct6kRXn2sh6X8Je19QZcLjbw304ws38fnuTNVxtqeNy
D1dcCvK0/mNgScDH7aqQx9zbo/QECjWY+rGpHzaC7sBed2Z7txo/dA+mdQkxr+y+Fs2v3i3YxB3c
iQXIQWhsRSPi1ofECxxGFq+4VB9DX9dE7WIctfTFAl1JoxayjxENjqkuL5QCb6lgxO2nZVIAkBkR
PqIwqHPsaBT8P0iqCPxId0Ig+MfkYwsp8ZluteQpLBdQNxlO0a/OCmVlKKRYfT7vGFU/cSa/0vkp
xGW15IgOOWS1zgguk5lh/OCDY1HW5ZF7xop5aGaToo2ro3VGUDK6thv+AA9ysmuRIq1vo3+y1Dbe
bH/K1NDhnuJiFAo2IjWoPToRwCzStltzuCExiAG2S+MXVUHxyDKDUnfA8Q1koA/AyUxwVDYLa8Dr
x7YBRwr9UhhRibgmyxFkrBkA9/dqceD1KIrdFpwfI19bkviDf1J3+cqDtcltRVdnbhYsXXNT7Kdj
yzvZhrFLHqVQjLSfoDREU+TOEJYqEDO3DnFogtQzWwV9lvaqofDwMfqX27+z+El9+5c5TCVyKnPE
P+UbI7ONyCpSczLQZ/AHy2mDIwuAiBdMfWMgv1+hjbkAisayiJ3CcWFGdWJebwBCWXl5y7Ydt0uQ
t/wnmWdCU+goYd1tfzfeXB1yEfguQlT550jbEs+4DebMoj9MWQl8sB7nMYj4b1sNcTvcisjDro5O
Lqq5D2OLGfSxBr6UUKvopXkQ66Pq4klt/JXF6YmuqFk7x6PRoOC3bS45woa1UW1Ji8OZ96ikF9tw
2Xdwmd/e4sHZz0g7K7o+f7b+hu3r+FD9Vjx9CaxWslWWmLRc/NMi/P7E/SYlOE9jnfRg2XTayBy2
n+orgkgSlGBHYCEP6hJ/XjaxvkOC9ev7nRB7JjH64A68WPmCGM5MakZatKkfEoJ35MiKDNG8J1gZ
Guhas6UybvcsM5ntamlmDPFw4/VWcI4SI9AaMMPXelBSi9kqj4HOlbjXClwDU9KeWAvuGJcIDcwf
8/3L+9QeAuWuLRY1UdOYcMI3ebZbmCnFGBRAAYg0e72Y8RQW53/mpP2MabPu6elRbL5WtWbaTmnq
BHRIrL8zU9d6TuAtMb5Rfmy6GX0/qDE6UBxBWXKWArCYM02qMaxCcpJL+YRX5vJP9mHFNMHmZVYC
O5FnITfPsEh9DlD1x8HAAuiWzWckfIKQgepLcqilqz7G8DYSCsyIEXlzq30b3Yar9Qk1/R3NWCNA
PTHeH1c+ccMb4fI209dsPACKx/YPsjEvdNUR7FJ/Yil3EoK36ruax0RlOEmMQe5sbygbaFuM6OR0
9tS1tLIY2abuCZRJVqvy3KXXXHeAhB5VFuxof0MIWBNWMIKSE/kYSSSbsC0cJoAamt8gFvoRc708
xuDoitE6a1YmaSSMSccRECH1GpFLb+UTBbdtS9dMcn4s9qZZNuAYuEHpI3wQ1lHak60Cje8/LBfK
BgLZukNrVOM0KLlLgUDfn2MoVrR3IFeIBxJCAMrcDibzJmrBM77rx0qqtCbqiVbyhgUF82ObCkJR
y5O4uWNG45pRBUY7LLjvsZ2JHSllwqT71JHQHzUbtVJIDxAGlw1Hv8ddoPiK66TAsMWYU0FE19pa
T1lrNNKbCw+cBhTpCo74IWD9zKWhJltand1NbzvCtS6Dplmknq0x+/LKO3Kn3NXU6XhOzIjOsHna
iUPfWDxcilw6Sp5/gaPHseDw6tOwzuCE2j9diEtf3uJ9EoGkdg8UlXcsZtVldEm259/LYmqEmcYS
vFUFoqUsjxAk8GF09w9wo1+WxXQNlKKQzM68IxKNhvOUnmUQ+LQw2NEsUhImz1xBc1/FFDKbEBKz
fDQT5GABskNHN5cDlvBO4L0qUWzj6QbsQzc2cDBvNg8472f43DjlQCSzfZUTrbYioMUNg6OWFWrk
dLj3+9mjOD2B3Xy0Jy53uz4806AtFSf9Dzz3vvEROJleOffDuzB0QKbp2xPCJE0DQ97WvJHAKafK
mqzIzi34prPFwoEjBDTph5EEw+cjdAl8+MRW3HN050p+UbgcXqmuL0ZsM+Ehkyt9HyRMAHEzzAM5
GR//q5HjzaVG0NGfM01zI0X+0vX95ORYFauDWSfhOZ2wlpxkbYu2rM3Ti2WH/J6qUayMlvpqFbVC
DmHJJDE1/Q3W9+DQme5SC+fcrHqF/XL43N+qdCIUYYQE6gJE6LCLL/3jJSW8U1Li/xYpb3Z0gg3i
MxWG4hTGlpgGUiDcntun0dL/AqMN9k7PRmWISe8jgvaGD7RBR/+xI39LGm7TW+mJKUM1SgPv826H
dqMS0mGa2LFuIRQOFN28GBNPYii+U/Et9RmGzQkSRIPvX407DMSjrAxeAGz6Lj73BMAinVcY2/YZ
Ymcu5LhhWWeZcJ72aYobk3ocIxSH8yvvhLUTOrmrPv5b8CJ9z2cHmjPogHFtF5eVq/UNduOXkcRx
adyOQ+BbQPISYL69sbZrKP7QHbrgL5NHEY+9f1RFqAyyldIezyHS8s5+QugZBzVXIaSV3gupCFRJ
aJXRIh2FovyJALTPL9Q1yVNYbjaKyJtNKl6yuPAJKqAwJUEVRaRpSOKWt/oSGfvjeZZY10M0YiH5
lOVYk31k0O4DUgtIXqIpzAaSPj4M9qmRVk1UnfW1qGJiUaRF6KrYKkXzawbs+nQx+gOnZGIJxB3p
uDukcsoxJ8SQhMTKYq7iwZAsnecQoVlM6So/VmfJ9YLE0837Ce3y46kw2avoTfz3dY0FJ8OciMD3
QUNyGo4kNy86guuQvMDJIC4N99nm2Y3L8tr1JvGwcUFDIKx8X120LYkU7Lb6lTdGIKzxeUWyfv3P
h9LkNV/NNxMJl66cqXkyCjdeqdYR9xr48rUNANaltlkS8h+kMeUnv5BdsqvuiS+k1eLKCOvcSXEp
lTZ8ZhKltSMsjop0OlAXsGStR9e76kZkCs18NQcd9rUR4oczu/OC82HKv5H45rI6Tf1PkcjsvaRB
/3JBr8JeS/YBx5GYyP0UpkgKA0SkboUbJ5QlZEuQ6lBJLmpmh366XPwWahHupoqXwTBQltAw9x61
CZcsbUvNCIyq73jzYH95v2w+mx5DWXOq4owYjkt4bkIZkCKdaC50ON69uayZ7yi+KOqFXIJ/m7og
S/hZGyByDfTSr+6ll06juTCa/mO7JZBZL1EW2B20LaMAwwondg7TD8B+eYd7ydVwiIubW/dA1lTL
GR07Jrg4DAWlO1CEc2OyAI3WxZx258shEgICJ2pOchNYmseqrnQEGaUB87bY9ykLQ4d16e0AeR6/
7ThEEOvGLaqYNjONOCp+rzSqnqtVg66YHWMemw0te6i+7lmmCcnHFzvckhyeMzObk6DDjwbNZlTh
TUjtgo9J368PNR3nN4F1TxQ/UQNCooMG7RJgZetBRnEz3G8cXjz2Q0ngpHSnCKceIoZrHUShd8BA
YHKOFZvcYq5CIvdBm8FP1xsWo951TO4QP1INBhACKxeoV5VcWXGK8x7GkApjJ8nYVVwql8RRTq+i
lS4ONXVlQ8pDepg66yXhxRxzqv9otOqGEEzeIRl4Rv3j90rP3YVqECu5lknBUVMqQdc8Z6Jy58us
WwZoErxYuXyTtc089eoU9t9pEqdK4Qrqdld+FpLmGrhE1Z6OG6w8ApuTxBTIakTTxXCQS9pxEd5M
DIis1JdaKOHjFfq+MJGPiccMlbBaqP/WPBo+g0Of8SfBmzAbcPmZOwotYb2+439FuSa5Q2025IaG
7X/OqufiQHpPXykHyp8omImQL6COzAQMUt/7cepCHA3Kc8Yx78zvch2Uur77qdFdgJIAYq7RLrcc
gSThnkQ4gn34sYMz26W0+DXpCEJ5jh9O0xwhk1iGXYi2R9RSS32i2TJQ9uJZRfgLChjf0dTJ6+k5
zjpJw6iN0IyyQYt0TK/kjr4pyqa9phef0FKEh3LxBt/gh1XGcFpsyRsqw6EFJUCbGTFMNFUiBg5s
KJH6FgkLDj5BDKNNoVgp5gQ0h3NClA1PTZvF4POIG+gi3KJJfwGY9YzDevQqZ/9GnXnqGgUNsVnA
5EfVz7+IsHuNwzWK6dDjMMwF8gImGyms+YnlFuozdvYxdBwxkx6HGenyUkt7lm8bCsRo9ZQ3m9W6
sQflok1inkmP65xZ20zEwft6/D7XOCF5jVAVUc0AVNjrOj96Ki8MH5BfBkFKst0UUDLyttomQ5ly
9ufDiMq+VJoXgH4Z0hcxIhXg7+oGNTwjB5BPXRe73B8G6YexkD7370AxRsSR7Cpv/St8cbKhf8dY
Ndb3bUAmElTLW5v4ZlwYrwWJHA9Ip8YSgu1//JcP8TS366FPjx2+4GIpxYJCyHn0FmQo5CWIqLbq
RkA0Ta7okOT+U0Q/ZIk4CVgLlJti34TaC2YmGy+n841FU5BggRNx7M5RJXXfWXpi4hf3zvQyRMK9
bZGHO/h6+88LElm/szIpTjobc+gzayXj6D6GQyEXShf3FHdOpESAqazooXtIze1UTaILv1PrQUf4
sHNUfNyvTohGZF2LzBvzt2uqHzIGYpv92C0afxZzp5Cq8Hpr9oorcPcO8u4alXF1DDATTnbjnDWs
paAN9GNWETlb3YYPUt2kS9xCF0nnty1nOT63UB0DxY8exroiQSUI4CY+b+yBFzgBLBgehHQu1NiR
9u0kt86cd07cmGU6L7JlYHMglFJjLzymBLAkE8mVIxVAVN2D6uFffT6FL9OncFyCYz8y3V08wPW9
339T5rk6xMol3gUZwW4S/hdB5xwSHmRsn0eZQG93OdQ10GGONbL+zX9DjvSG0iRhfvSKo+gM4Rzi
bG0CKvg3H1vliHQBBhBImPA+9xlJBrS/+XiehWLOIoA9lOCbxPCv1Sci/oOxQm/NNNbGMKz/vRpV
/PWzRF9/SLVsyYlVAMhjOn0FEW5MHhpMCUWFsbXw53qtOXkPG7u20wAe1yXDTsCMekDv/i/4VXYu
iuDW2rYQcLseiYIMMSn+/E0MFlYMRmIp7hykG/eePft31ShY7D6xZeYMpyOVjyMcYWaFcX/hXA3z
tPbq3BWAY3UpZCYz9lnFMUbxPbhR1TomMov2XzoseU3i3jyMlcr1CMlTrNd4zOzd9e8/j2Rpe4aA
6JfrbeHZjuft2sBzUpgWjQ713H29DfLRuoyPaXozlka2n4PpfIDVduqpefp6s/Wxw0CiWU4dyjfL
/n0Uwa0u0UXYFobcF/bo02DS0i+Lr2bi7YSvGmdg9Z93qIOQNrgvV70F376tlbFkkdGMUwkFuB1d
BSHsBhxUSWKOorzRnpCPIUbJRElJN9ILjPounLBcy2HxzVaz+xK+k7Cqjwoi9Wgovv94iZVejquV
2Q8M1DkAf2W/8ezRtpBoWxkRfs0/pRmsnugxqTAYYJ/rI11aJ49VU0He6JHbEgNbzYS823/zbdaT
QFGGZMHG3RnTkYnsOJICjooDIwx7DwD1Fs+DMoLolU0dDpeLzZ8v85x8fNcDjHB9nqRIQt4s+4gL
6Odpf8DUR2Wiq8helTk1dLDtCP08Bdtdh3/QG9pUvlsYOOaVPK/3S/ECLFk5p43iiWYX/Ij2tSMf
GNZTUkjhPJnGMfvSYTY+ucyMcwoAHUJp0RQunNsYHMclvPUP6xIjGfWNdRctBX0BmvjoRJgVp5yT
oVRkUrjiL2E3ltjHP3zyi2lN419fnmw3I2fL3bHGhscLxp/d/Df46h7qQMQYfkMEGQrPyGIE7X25
xslvMfEhZ/YvSbLVHImWDI23ZYahgSS05YdiTh7UmzdGnbIn3eTfTKOyd8oSjd/IZIFba9CKfMeZ
GXvyfPEVPlBBVfI/eM86s9KWOEtVID+A1UlIllWZqyAZqv26WMjoZRbeS+ARetvh12iIbJjRQcah
lql+0GUNP8SyBBt3aaDqr75kJnRrwksxOSxtfzSUu9CIjv6Sun8PzUlS6hm/pkGaPxd9M1OPYCWj
rKrVmPBwRLoAVS94cfN7SgHWrNr8kW6aeSuAWXZpTa22JvdjDe1ggDJ/V9RbAQh19gRqNls65LLH
J1JImB6F+Y9rDHJjnprIq3SY23poGmwHjoZlhwTvR4W9vv9QbGkNgo3LjcIWvcSjmGzyZHzN/Hhd
XxjtdzZRhX5/x2jNl/yBUGapL/u/0dUCb4MiG5Niz/OOgmJIKWjs4NAniz55Gp/6kabvUa314hpA
MHroUFVzeZfIJUxhGiVnpKGW/Chb/u9y/w/Yz4QLK91T6h+4Rl3plnnFWqQZyRAHkny5IDgv571e
xV+lQ8AzS6gNuFM6JgCnFLCIiefw+APm0mhXuby/GN6ezIbRp+4xcSexNZrL7G2L17bEHTlWPC47
2YRcTOZeXfk7joCU0M8FgtdV+Pat5ONcYARCTLtrsaR+rVnlOdalF+ljrPys5TjeZZRpQ3JncGRq
WDeJ+/5v9+7MmmRzf/gYsJuzM98uvpVlKLEFuiGTotUtvumjJY70i8C62IMmm+mqrXlQIBmM8HuQ
YAlASVR+2DC1jdumF7xPFKXdwCLL9c7i2GXU3w2ptkbUM2Mfx0e3JMDaKs37AjOhQqpR7vnpCrTi
hWNh1GgjrsMXscVZoA36TB06FGL+YumSMJauvFKt3Qpak0sZhAwVDFLEAz/FAur++Ge6yo1KT5zc
+pobsiT1XcYCQT5lj7CyWK4p+yRik3Zi/eCd874rOoA8wWhr/OnNgiZJrME5L9auFwuwqCoviPvt
t9oV3s06o3MTcFIcHSHznic6pE2LlEV8M41+t1Mrl8+A5xhjBKx7ZWM16p5GiK1YelxpQVO4Eymt
lCUaPV5agNwJGmxca1uoWyAbd6nUNmMFpoD5bmz7SVkb8KEi5OkyG3NRpp8cjXZd7uVHQ3fewxqf
qxI/5y7pL+yPCUAXtD7AI5AySdDaSxtn+UNyOqoPyv0fKApliXmvUgNiJuXUvPE95cLi6qo4kmO5
sAZ4obEoHk4F3joynxPoBGCD8XdI4itc12IDnH2OTj5hlM5zftDfruI2WfEk/eeZx6DHaqtcJ8jn
WldE74ZHzdesiEZpb3M9oN2lkb1D3X8H+ANoTDYcqlqHMeRlyrJUlQ0VqneBJD+JGfzHOJDm/qg7
8eNjIheT/jUAEQBxlKkh9v/N6/ediNvIhQYG1UQaFx1QJdtYwp5J9yvZaPeWp/b80sauK2rB8E60
gQnkrV0lWNpEA9whMYmhh4hiLQJT49AqNk+zxKRqTKGh/9NsnMDJCPTyTDmkowYaP0YWFAuYeMAs
jfuTN/lqtWlcfEUGjd6hwM4Ynrq7LGZSroOQ8DP9w+HB1lS3oJ/DiDSglhDvraHJWHTmkCEX8bVi
511AtBnDMtlSrUQ80l4lkfdHrvyi/STSxMCgP2cJYukplvIZMJT3OYJhb6GtP3v4iT8C5aA4KPAj
la+SNQQ/orDEovpRPDiIssFvmx3ZJWYTmpliW9QWqXE2pmD8LInHg9/xTvQ8AkSwJyFdJxc3Dw6t
7Wo5Zcdx9NNrTsvkUVE+wgh0n1MO02JPAun5TVlfnWx1KWytuiXRzNQMs34ZGr20WMq7iMIqp7QO
R1SO0On+hoRJhAti/dvhF1DVXyy+uRvpo+CHH8MQXmMXblL1VFctXkem5xKClyf0pfIo+d1MBIPR
+iqi21lEUWBH0PwOBM0GYDxezq1aSAnwDPVL0Usl7VmjTqw591IH9IhMdPd8nnUMEB7lh9hVvCCp
iex3c95LVvlVxW0YpHbNcd4L1iKwTrs3AQlejneQRv2WjRCzajhJZRw6tSnwylNs5rqGgrQXJR2H
qTa1AeYlxblGb85RKwcr+/D8NVMTSzBCrg8nkIeuvRy+Np5CpPRXxYEyWfu6W9lkuqYn4t667TPx
Yjrl87Zft4DkfqKReJ44ujVRWCrz7QMiFej+SobjbmarAKk8cXRkQOT2646vGVCLHLpC49grz1TS
NHHm4UCJZZCKOS2jogyEeHqze9wvIhvnSm/UOM1LQl2pH5XZ0iGU1gZfAVTQJzFK6s+dfs0ImIbi
vIcR2U2anaMBpHZS7dDVo2WHHTevVkIdoib1VhQ5skKnsOTM+UtkqkNPbXNRbWNUzhdH1vRQ4IoD
dvdeeP0nA56tnCAx2Ikb60IwlDHcvWmUCyrR7IJ5nvNxaTHBX1/MOPhsA3aEJ6FNbpnsrJlOpDFd
qQQxmhmVHt9Q/+9rpZfPgCVUcmwKLkNUxfI4CkxrHo2giOkUVCCmPfikD8ImUi02WfEAJ9Lo0xvM
lPVihuIJWiqq4i6SRKXX8VCOcaG1IyUvAiGyCGNbSyGNU7KFhT/Ccl5Y3hHQhI2amSuMAu0JmVyx
ZXCdh31QJuVuvRcoTlIqvJQ2EigloKozsK6f0YTMIf40LDth7jZoPX+ChQ67NScLbSNgZx7RDV+t
9C51nqNxZe4QzMtdRE0OXAiUAbaeQwsdfr89orTBMhOC+VAG/SLOXp2RdWE2pXiUa1BAZxa8gMjq
LQOjNdiVHU7cQI2Vdy+68dT+ACSUyA+2QBfRgb678LUqs67ZrwX8dptHtTuq2AbU3wok1rGrqOZs
5MYl1O2NmR3e4MxrZuYzH+KJpaz/KxFR0FUzXE/NvzV71kwjpiNKCk9v2WPd16oEJWDMJyfUcDcB
BWaMlGsfJ0uK69M5/XprbLWTcoNLoaAZYQ6qUF4QvtJ5BVra7TFPUbwyyFFmGhuSX0V1DFv6Onpk
5mf4kXCNddkeYo2+Vq5SeqmvgSdMa5Apnkqf42wdrBEi5dSpm+MNQ+SyiD+Xym/Mx55NEBKVdapU
993N6Ks/yo2jh964kY2WFYX+UWYe1aY39aZGparafbICZCAERrsgcGn3VIYCCPFKgCU4ueDpT2/W
1wN5aNxiz9dpu2vxLOEMW4UnhmNcqxaRRkGcwf5oC9VBZXMxmSbbgmvroGoSISeOC9VoRac3nCxC
uSY+gXpeAFnJtcLwqT8IjQMDIaPu5y807zgCeDt80oYcnaFlfZw9OhYmA8unvpnRxLd5yVrGB6Tt
P6f6aVNIaXrcWqotcV8wbKBf8b8zl5170l6Tpi8gd9LGWTwfdoPCZPHjYvghCAY0Lf6i/GK4os6E
+Mgqtp4MwURX15kMU7Tqp8aldNkxPi/OYHsRtINOP7pc8ITlboZa4/YR/fvgNfAz7vfeWg/nAkRk
XUK/VD21I7Pbp7/7W+/KG6CQA9UuhHQ8F6BFgYaNky94BGsNfMN2Lmwl+xIGwCdcGk7svCfW6iDT
Ux3TJ9oQciynLdhs45cCKtgfKAcIb2W2HVs8bNxluWbUiS9c1qAdIMlmWr8gzEptDeA1Dd8DAENh
EltVqHpYFbt5KSZwyhmoQsHIFQLTCLxL04iTMehQrsEnB95Cm+XUvOGGRGMFaiF+mLpDiVPKYIeE
DxXuUeRv2A8oWcEIswJ3SPYk3/G6PGZdgPYml3oHOUDreRxUIZPbFk3a/VmQZ73YMgpczI7iXfvK
vgiGmyjbmGYa/i1EEguLH3uZGp5w//F/u7DdqZ3jBkbt1BBu9SHnJ3OaY2f8ybMtRwXTFznCJFq8
4FQqCge1Em/L4dmA8uS00ue/y5EfTPPYQAYIfAd2OfLCdMW5zwRZvZxexjeRrBftwM/9vWGyAg//
/u1TC/zNpzQGRYF9Y8rpALF0XC5m7W3itYILO6IsBQneTDCk5MTnBXsCr5hJyDaZJ2IIMuhz8XOG
V1/Y29/Vqs/cio8KyLb+FZheETCGQnwP+empIn6/XrkIe+65yffG6ynMDHlUV9yUYBiBf95v3/3D
eS7hgdiOOy5axvHO2f5FLZ1/X49Avfs1rCyMi09mgu/zVBTWsstbRRupJ6JykX9mngLYwdXthV3G
XA3yqBDNA51+EvRX6HDxdYiAlXVJDXSThAE5s40uxARjxPDv6HwOOQtZ6ABAOPdNh6XrskNhmUpf
+He6XdV+/i/6B3whOq+6S0NKinUKTnlHPoCJnvWxN8hxk0vwMR/qCj5ia0yqrwvO3E8wdVUTMzYL
//5bN0fM642e2QWJUyGvat2Y3LI/FdsV/ujK0TCfFtvDnRiOyBntU21fwxNM1NjjyOmqN510RMnb
Kr37PEDGLg3TuQhjp9zdXD+nAN1vj0VzTz0SmdotNvnVAwEmZ9+9BxkByilRJQNb+Dyad+2i9r/c
brd+XsKHfRoJW04FU63huAIK2RsOrGATv6+ltbuVnLHc/ykCV9tRa4tT2/1FZmcHbqM+E66Kg4oN
/Hkc8AmxDRHl68UUtU7HkyOt+jgaBnAZS595QXw8adN1IZID/VqwG8yyBQ72o/EH51nWp2Lm2BtC
q1y3b1GSbT9VMlpedev2LpNVYX89MZSWCHKxrcXgEUlM/c0Tu+xvHdAg/CmEFsomjRN+LN5xG4sP
+4Bp9CYcCcWcrS37Bj4DrZwj5nnEWlOlscA/8RXzDT5DPJZ9CrmAVvbhSVTZ0yBsBTZilpjfrhDT
/eI/FkAaGilyNylcfhAzlBuhXzsAsBablI2qlpCWjg27xFg7alP+bE1mxjQVnKX+Qw8ToeSV/n5h
jlUB+YN6DG23y5FaWdaFiaM2wtxj4UqV6dS+FcY1skWS9X08ta+B9BkkJIA5A7NcaleSDtrPzGti
64p9jdbIWPuCZT1jJ2UFAGhpJ0yAVTtMSpDjDQ6RHEuvVTqQ+L8RLLHUXutbrjYDbDkcxOFAsBZG
xq8xTp6asq4p+E066DT1djjy7qsOJvo9JiuRPijpruO3rUSxBPpMmQFnVGzcJ31UqWb1tGoVW9/w
+rQibb4tbOWhw/FlD8JZSU3ETyuesKQN37xZrwAWrwulRfLWPwgRoFyfTaTO8tghSCsNaedxJl0i
Gl2ROWu2c5W1LVfuLk9Oevf2NDzSY8S+EerlkfYdITufAU/Z/15HXoPgb5Sj50VzfDZ3B2hwLNsK
TdFTkhH4kejLWPgfOG4uBerzuwmjxvHlVMByB4UjOf1QUInE2ggyCWNdwwWonVux3kFzVABhX6g/
41cUCYSb4gkjTnR/hX1jXDAmkbYaB2V3CYJLK1NdZFcrYaqHlA9bJPUod2TtXABc2QfhtXdq945i
biLR6yyow81YJHG3AK37rhKyhMMBehe8Y+fkLmSABtCgq4XhG/mgsd+GcsDoq/3OPakDSMRUwfrq
Z70vwP3VaP6cE7HixCGLg3xQW0i1M3VbLkMKPt1NJD3VrGZ+/qo6YxLmOHfRXk9uqdNzo8KGfSgZ
VCe7ACaMbd7OFRHr1fIii8vMFZkJOP295mQpozr+GPVMtI81wnOWdeOx2J66hYVijwkvCimlcNsL
qNws53A39XyZw9qc98YIcqNjPTh/EvYjg3syyASwaLETyt4A9SfxhreUKZqoWAqEUlqNldnOLLfU
8YGa1sE1m2tpbo1tBYJj2S72FxfcQgRvNuEm6qPZPjOFrFzghu+bUFcGjsq1/xCZxAePhwCzrau3
lwWYq2oU/hA6rLKWmp6ie+ByAD6kYi9zE1Jy7WOlRVjAAIoibcbRccBWRfmt7Kd+W1nUAx5cwZP2
SiLO1FL8bTj7l/Fqm3jFOlf9/NzJijj7iao30hytOaAWmgsI8MH2MOD0LL4ZmowV0JHseZfXIQtn
yRafUPdydcIZLiOk7sOkczC0MX1nC3rjvfxpSLkF/RngqGvCb04VrvXeEn7SXtr65OI/qLVpNeMK
M1S2zEBHMXEHeCatSbatOuj/xpxEbBrGm7p8G2o6BlkHr3sL093mGxFGgEYAs2fsl7abCr8cixlj
vI17fYCbyIy/AUu0KadPrl0167VHFo5vKi2HgiBZNs2CMQNLfrQ971MLU/xW3MtW6Okg8hhvS/Sh
1ycabyDuhx3R9Xg058K4aPYI+KYe2W/28W8ZdLac4KZ7IfylOJahEkwDYC/amL0/r1YU7wAz1mBK
3vcxZw/0/UUII1RWYRyPMI7454jT9nG5TFXa9HZd/VfUX72o2YlZAG74qb2Elm1XaWG3X77nZVaI
FN/uz8Yc40AFUsZYDHEZWAxuWIizqHqIvUsg7YfopMCy8L9k7Uj1suMgDWdWKuuWATWoEEn6aELp
QJmKb573irtLH5uPx+reqWnpFAMRP6vKnBghidoMcKB7H9vMZ4WlX+AfEdHabPzEx4pB3cgcfALT
AriBDBC/+ZdZ2RQ68RdqgSeVq4wRftmO1aU2kKt6+mQPfs9avO7x9RShmLvmpp4ylZUnAqND4tCz
l9Mkbh4Y0hlQtzhQQ99mmTRQUbCZTAXBWb/MzpBccoYhg9OXTd8BWiE9SiHLGPy2ySWd4pUH685h
uVB604DFnDiSW1XQh6D7BMe6v1eTdbrW5aw77KDLmeOb6MEydnxgZw0Uchc/n2k1rThlXa7CTMsB
5m6nVcpKvo7H5PgJc84RkrGXMC67lCgr4ZlLQSSTHNSw1R6CpOtV4lNzvTGgsCs/71cHnA9mwaqb
G0FkFgNveGTSKYIUBtL8z9v1x40BobVWclHYHw73QD3cRx5/j7zhY1MXa5HyBM+9X8DQyhXxO/ba
1TXlVwA8Un43ixZ2GpFoAWq9A9pHDZHGfbkNAdipfC79swHIc1UTN/SfDYO50ltMVTFFGms3U3iC
M0DvkhmZMjQvo33Nk6yvdBS0Hyv71LzG84M4vQt+ZT046vTpk6lfdv5GWC2j+lvtKKA0dthwDJxH
IP0J1hyFi6IfJCCau8e/rCzNJpbhTlN7ewEJDOUnl1nfaUVt9vaD3lwctFVQymSzyrbSbxUbNL5T
eR+P9ypAJfbI69Hm0YeuEaxfmM7vymTg4s56aBwjgnUl4QPMJmXuBpb+ESXbHONHgRmcSBH6P7ie
Mcjhj02YloS+1xVgkeYzKtCOXYGWNDf69luiMtdCD0MRDwgmJGc/cWMJZ1tgVhCIagLN9JVkhzpg
UDKboRVnKQ0evTopqe2xsQd7LaYRuxbS51PvPFWJoSJsJHPZDVtChX1NsR30+sdGfhqOHbro2Kao
hw+VXCSlNCfRxILOJmQ0z7a5T//3kznHgwzDIVWaCzfuKxJ7nm3DBLa1K+EmplrGsDcIEywxP1ZN
k2lAQyDEaRb/fIaIK4NptgkCgEsZLnqVQIoA1IcmAXSrD31FgOcoXMsdllcZeAEQNvYCJntFTkUP
8K4OySBlWonBH3q507AKofV8eHl8dIh0J3Wq1FLnslqEjjmMDPN88Oa1I3DlE0LDtHswKDv664VC
FENkcm/bTiZ5Xwo5iRt00Z/XSf1h6qfzhsDo1yieCinVjOlEkZsRuDxQFsnmxXBphDZVhaLACHk0
CaD0IJYX/oIsisZr+V2qoMgZl1DAIDucd5D1GPp+6KZvQqJHPeKBbjLUa4IoNB2QIsHpiMJzGJUy
ItVr/vmHbpmilDKx5538X0sA2Pu/2cC2fXoKojRVZCv79xFsEBIWdfHCZzJvOELiAssGzWGbD5Sr
2cnt3Gi12VZaCBgYBgPJH6/ZGXWWTgezAZBiPdg6W0ZuELf4meAhXYuJQPODHTzHO0X45B0d7E1m
HHW+JskWvx9j/+vXlY3dP2+wh4i5Tm+ACM8VDEhwQcWMr/C/leQqqu+5QJWQjpN13Gqs5yqIT1MF
TCe8SmgTFCnPe8vdXITpkfyn9J8ogYsYwd1bNHEZhModLafp5DBdWbIp+7mOp0+SIQ3+S/xIq4O6
b0iI6QhgOonFw0582qTYLDHbkwlnpT7PyefmavcMxz7N7Pm32KkTdl7caNUHRvVLbsJCFSwpi80V
91c+DeIlwwsaSJ1AgkHgaxnk75yuMHXt1OFpXGqK0EBMsc6KWI2xsPYPUe3wCwbbhmKGjRNDTl/j
kSX1HMQ5Ddx1WrpXYViOqjlSVkxUUu+O1ovbwHSOVOe3PwAWnGT0C55yPpLAThPIEJexmT1Pt8Sn
jCVOPmdICJM5T7oFXx2o9DZ5T2tUdXy0BpXp8ZhNws9O1pZcIhUh910t1hyN0V7ecm5vrHlBHWB9
88ZqvuoTN8v4xIkr1qN1TVUszEKrbgU8FHt0o7C7mBc+Ex1kGBCYPYkKlljvEiTKURguseExlxGL
8GqJ8SZifNl/HcS07VyYh6P0TpT8Hip6TtloHD7siOB4YD2NsDCSaxqg/+3oO70c2kJk44mvKRSQ
u7a9A4ZsHO5tmd45e9+SjHKhA3rkUXtnGQ67yVS78gsF27hlCM+APv3Jl4uvpSncbnns6xyaUmXG
dxNunO3+gTloyVqEaGwNkrETCSF41sxYxxitWy8r4ewDDraewmK8rQlRcaXMlqiItKCjG8Q4iU2L
qEPe0ULaLbsfcjwmOPGV/HD5rPKoU9od1AL4vfP+kwWKfr2xJOOT01UXiq5sIptCq4Db7omFF7aL
Iv9dynSHCNNI3kgaoQIbQKaK81zjKNuAfG7F4eG/qct1tNi8iJ360EtUp6WBSpA86OuEGxwiAHbB
ViJdsRGb6lf4qWX4b8wJ1taFKRZbOBNdalRSEbnPiYdp7osH5eBYwslUdsYXQHqwXu2q6kb+07Rr
bJiWyEuwg+UNOrXPQAKrXd94Vr5QEXqPd8P4IR7aAfmnIQBlUmC6miycyxBVLnsAuL4x5K6igpIZ
kLIOENLEJ5ms+uzzGaqQPB/z9A6QhUUofkdXfvdAeKt8QbrTBb0RIK/1sTEkRwkAJp4LnTA5dNzT
0ygqEDhoG/+ZA9v3LW5fF2uSUbNYyVoLlInPeCj/kbvkmAYCjSoFMUewgJtTa1tq2G3GU3ByDHrO
j06xca4/cHmiMP0twFSIIJWt/I0O6lMXVRzKZRzt0Pd1jlinVhWQGnyJBjp4svH5tf7QWbT7wFHH
gi/3ZS/tFu/WDtf3/8l1Vj6Qb0HI+/ttt5BAM8CBNyX8MyWjbt9wqAu+0t30f/RVavheft9aqsep
Y66s/XBCz1QKvI9jT8sWnG9PBmN+X1u8ge/tBXcJ1sLqKj5+RfzBriyMeGKTXhT/LGxZ+UIzsI33
S4hm5gY4sLckv1QmaWces+hpDsfYuwYKpD/NDhXHaUQFkAPtzz7drEIqrgK7MrjoViLNFAV85Efe
n5ihOmdiFczCrjP3BfjIHG9r3FtN4CbPeKHEoZkmXPsEVa82fIIYl2wLH7gzbOjE1ku+zVVbVWHO
of0KDwoYkLIt91zBjUufyt9TwNUI0OaSVrBoTwMTM8hRWO05bZxOry3sZEpgFiBsMHhD6+p+3OzF
yPz4iqhbL/aCMVZcs9AFEonXznxbPQaMsp5h5xqYeszZtxXK5cC7LqVuCsoY2URc2rhsR/A5C/Hx
Auu8JF4tLvy9vpmxIDH9e8iidrNGdKznAK7Hi/pncVkGDTGcZzz1GahsEdhLGFFdk3FXWh2VUrEl
QQOfC0pWO74xaRHknVzPsyyhu5CJIq4rpGqGhAPHqmCkJX14GyGhrKjxOSyTp7ekd3HnTWXV89Bp
zEac+P8cGaL1Y7FKHPvvr9y1ZjzeRxzlpZRtV1UkFyvZQdlRsS2DqH1OXVk9mnqGGddWMC5mEhYg
fUNCiOSFkbipPoQBj1Smvmla6K34UwIMnX61iZuLG2yPm8wQ4d6NVkEGMVWCGy5rSS8f4kXVzwEo
dSdmSUGfMrDnNNIeYSlS+Q2q1WBkolDX1a49UUxUfBj3YLfYuI3AgciI+UBcdRYhPWqbgi2p5wLj
M24/wa7ovLDKZaQPkHHISPABlDO3S41mQOvcPd7oTDNEfettslPK4LO0BfpEjSemWbwtDD2Vlhm2
Mtl9wvdzTstTtN+MwJwbmr6hBmY7PSBnd/Xlb2EhSt4UgGm/r7iPASg6GABusuKimR1uJc06rv++
Opf2lUuFMqS1QQ8udNLE27GNhPbxGYnEgFoDybi6zj2yVIAyAfQbUYOwp68sl7dk1b7ESoYigE2B
nlzCIDjkBeL0I9x7/LqytEyeXS8v8Vv45ZcsGrMbzQ9QwnVCNB54DKUqHT3lw030r4V2+LzSEVSN
a1hqqXU6SG25r1S55SSqH3KEiOeYKjD+IasHa+JHoQDUJ5UXpcqJoR8DqjHTT7sbTDCQG/YzGKdf
JTtOzLPTZEqljBpY7Po9CEflLFbc3ADzEJZWHGrKMejpIexPGu8/KqzJoFBKKyUpKT2dT87EkqMZ
t/KJ51v9XfaBY5fJF++GeaczO/FvDkxDD4Ap79PYPzRqn/j8r9tuItGjmBVG7gln3rKyLtkKFlJX
1XzU3ZO7YU0ZuMsStq6Tj6rBzoTt5HLuxEfdvTIsR32LnVL5pKwl8+5Xes0nXwohnl2vIG9ighZK
/0gRuioNmKS+0wCsAF5O1t5/7GKu8HFXhONQgBn0XT/7K61bEcBvDL+vpVlxBlCXv5Yoe2O9XwmK
AIe5jEEPwKUJsvtMkA1/C441wHfKhvC4Kv6jhDp3NBBRFH8Y6bzD/vPaEXk4XIX6YyyotAZPypK+
a+wpGafdeF6/Z7czBPaTdmkHazqlwT9k2pswXyOXadxeGtbrG4KmQSFrPLuVhxMkw2kRGE0IuY3W
S6z14i0aLpl/HjTbU8D26hIf+0LEWHiur62rIuqwpio1tfyCAi9Aek1lYX5fg3yRAiTpWrczXBFs
0ynqrG1nGnHcN55rh2KT5zIAe2pC8oAga739H724SwXxGpLhd8qHG52273GtEf5fiij+9v2FGv0E
wst1oA6d6ztfcEp7ilqK1tzmp/J1y5qvzdK4Nf0gW0Ak+ddpJ91IfQ7GcfS6vchby+SS/v+qsUuW
GKX2ufXA2ImkfpgEDltko4czRQPdZe5FxrPRC+UQxHuo6D92J0skm7yHULrAujl0VpihLmxEBvUo
PipNU32/fOZnA7oQelWB3arShnnMb6RtzUlAK9CESpVtH1ZmeSIQmYkMDxhX2PIStEGKug4/FoED
j2NXCygZI1GV0cPCxxmKRZ2iTYX91kavfcVwVAADkb0UYobYWeXQv5d29Da8qLPBGFZQ02bJNSix
ItwMn82FrRPAzEN4qsPnyHX6SozlqZF6k8ErBFJrdvl2YfMuJK83ORuLhVCSpyMsG1pme/a01h9i
GS+BeOHsD811ph4PZdIe2s76f0k7Pw86pHN77QRG0cC5oE6f7ogHF1mSG2jgdhA2k7Fppa1rVT0q
luRoi6SZSvHaCasYimG4YwPTU+WYRe489egDN9h14zd44tNTzpHioeUlxfADgNibOeUqQUrPsaNw
vCeTYeXZ7jiAi9u5zcF4ir+A92BW3r3Q42/potEBdduO6/REig5qKQyYqTVh6HJe/08Z9MIfuwaW
0VHN9bNBMujYcs1gNWmz3/BiVWDLZOkV/b3PYRWJ6iJsv/OdIVDqJSJPpiTANJkzglyOgi23zlDp
fN7QPGnYjYLMHCkEH6DK/H+qlhBzw5kK9QYE+ZTbE8vUp0vrSNv1mmfly5OgOOP41GYb2X9LfLAz
9zmU/5RwSZtnc0K9vLQY8maEEpvRFysVMWD7dq0koi4NvsdI2mA8T7SRRUX0zshb7fu6Uaiswumh
nXE+OK3sAf8CcmgBikEos1qRvZCFvh0qaBcrBiJX9PcOfjQyywO3i3tOg+ggbrinnHbULrsP3FnD
jyJBnwX2MfL0NhlEzuxH24FThRdt2VHfL8ODbWiJM37sWjysIxkhFnsokmH+Wle57acVxc1eTOcO
5yhinDzdHasR7Gocsyy5cPNZSvqaMAhvQu50soRqluqeb8J9MrlH4Zfa4+uhDaBeBSO7JwPU+I0q
HHyd/niHyZ1oOf4XZ3y+t2gzjR7rp+nY4rB64JlDwTbLxR6psOSGpFlxvWHnt0UyvG+y5DEY3UEY
+SAO2Ula9910eu/HYRJgnlSWeM4SlzBDqph3o5sHuzeiQmaZ3t4kGzqM+UuPwStS64KGohe6EXZN
Nlk1f5PlhG0FcTc7YjUqNMg2xA0NusA/YAgu+/czDTv8xn3DCIkv+vmaidgFaIXI0SjiGLFt9fTC
Wn4r/0wSG2a2LGa7HQz0jRzmVoUlle/uQIaIoW+GHLItMDKlYXkIzlyYBkO8OP1Tuai3dAhqsre6
XRG1ON1yB0esDNg72OzqU9JkedmfgFWT52kGLfZJSp+Hj41ATJfQAtcCy1OYPKDHYpNMP4CAYvYS
B8zrMx7wR1F7rJ/aQStHpSrSvCzH/GzSevLK08f9cJTdJmYRzw2+Obzf8R3+Uha32XXIyJN8OC80
iVQrh6gJlPfv/+CmdptX4zHF/JxQ8jRIQF0eOu4sAE3rGoGixO0DjpD6csir02SEo0vsnqYWInJ4
DJDlN2W1sLFnmTIe4eTlrtjCjTgt5Q0s7NE4WtS4AsSI18Joz06Tek7D3s6yojBa4vlTtbCJD5qP
HI1cxdVA57dkxCdXy2RGxpmvDr4pFvx0tWTpizqKVTyGUM765T//RsE1bgCbvzPD0b6Fqzu1F8Ez
e8HcpB8AMe2Le9PZBqTfchsFgryJkbSlJbdnWAe9+1q15/g5dnvzPCY/QNF56PFQ3XOUUb3BuKC0
fWm9BUIXw3ZQc24NG6VCMCG0VV4diQR0bxStVesKUkj0erIVJQWojRUvXpC0+rUhBl9WVx2BR4Qo
B1iEgP6K6d512ZioqYLoFcUXwLy7IqvsvhswTe/zrSzg7W3BPGV3tyByWM4FM+ixQuzS86jUItJx
A9ak0v/l+zAUEQ+U+vrhBxDViVCpWwI54OsPU5y/23RTJqKFWi5c+9Fq2YsEkezCVkSRG7c4sofs
+BE+CLmRoRAger/y4mXXeg/6VUsHzwQGAOtqJ8GzfOiTJxk6dtHnXKW5RRJ7pzqmhi4U4ZgRw8UZ
LzLYYJvbww09wWTTZHOUHTEYPSSCEfM55vIP4MolEEZXNbUXb+71QKS0NN9hGQlkU8ypiRU4GMRE
X0JwJ0iDFUEfXxH5wNZyrubp6tMAJVWHzTaXSIvwDoE0RDk7cTy0yQkOjwPNtaQwQcCn+0vpupIm
/25jNJUz0M1v0dv0l7dW8kSIK2YVvdcMSfH+VCax3Y1KCavQr6E4uKthr5DbR/6EcR59oYGlX9bU
cpIaQdKj02cQWjAOXae2TvZT/0+lUAkraKMLXnLEv3n2+puMXrqv2d+6z1TXAVkvypI5NO8ugaMJ
VT1Bam+YREqEmzwFb70Uc4LN78VKbitTNT5Nm0kGP9/ORF5B1/OW5k+5zIM/9nzn1x1f3dw1X5/O
rqqRam+YX2pWBjpMO6qc2JAA9kxq5ZvZiy2qxAPjbgZ2F84EYReGX+WRQ5DwySjduHkdxlKmIpHK
+s1JgWmR6FhFqd21jZ84nJK2WPLfXhAsxc9PIS9yEWfTljNldIY2IMhwnUYfhmfoUhOyR/oCl1B5
/bE24laEw5LxeL6wywtV/zzd8cprliOBFDlWQ2iBViQ/mBwd5QUHn08a5KkPBOOqCNZo+VZQELo+
AsQpUlF7GR8geJAzPXgn/4SCyg91231RHX2laM3zsVGzVcAHKxVocKwhv+CBlZkkETc9ir9ciOFC
SSS+QrtYgSXRjJWqEPZfLBSqPoQHxJLpfWlMkUgXffYu+hQzTbVdPbC8u0fCn7M+YU5uGq7GTTRk
Z66Ow/t3D13i6HgZIjMaUXUZZBPrxxikvt/XaAahlq8WnQY/JfSLFbEM+Pk6nXrSzTDYwS2bf95/
5BJSFNr7QyR5w2HE34Zb4kza2Lebif4oX4S9HMWAmLHYKs39JQyfwWbLDEYvEUOWApqUzh7cAMg2
OI2Vc/LLCKQowIaLuIY/2sO/WBc6oOradyOkeMvHfhVF+46pKZsWYal9IOP0BcWQuf7XLIIqvAES
5XVw/KXdNeQpdem7J17ANVIZg9SqjgsT1kncWlZ2eD4ObQPq8yRBd2f4+IKgyzSMjwxfiXfAvSu6
Odm5RTNzrmQZalLn+DmXNsyxJ+bEdZegHdjoo3EqrsQ9T7sl2VnOaplDnKuSZJoPHijJmSpJCYAO
GS6OccFEZrP9HobVOHWEmy5xvi7aPBSuAgGtaBp5/l+iHITTWoBReIRjd+U6c4yN+E0choH2StBW
ngZgI49531YAdTfJOmR3m6J0K8WAWiSYzdBbTauuX+62A1ofyzBaKmKOi+8N+K3r0RpKSiMo1DZI
9DWrRd2b7YAR4ohMO/2pm78tShKp7PDnyKvfGV8o3+dMGN5fxyqp0lYhDRuH0Yc4L0QrXidfM/Ym
3KSxEBhNN9oV7xBzExElXvy1D+61fjT0f6zI1ByNfJZsJ1EREDEm8iOrwRjdKL6MP5lpNiLmD2C/
usBg3z05ea15UtGkmiIasFjWNa2YwHO6jCW6PfZtNiK1nQR5Ntnu1wGCK4XQVXiHLYD87QUNDEgo
JHcfAGAKyAHDOb8S/nCyyhBrqvzYXc3NC+N4da9i/QQsMv4Fk4jQWAWgvugwqXEGCDwFJdYWxwj7
ZmoZBkbjQ+mdUeqk1Vvn3DuIaAi1bpKQEEULSFvQPuHRBrpG0uR3SN51FS1JeX7DmAVVy5RKNJJG
1Xo0+UTqD6q52r6wTR+ER5Yh+7cbVnpUxK4qhb0YPThZA5umentJR2N2Y0+7RhSbWmGQCYU150+o
SF0MWcadQ5M0zTmHlBHgfbgBxCScbcwplgGC+MO8AxnoeCUw3W50D1fqrzM7eXcjDPrsZ2pps8Xb
OVGXQqT6hOcq/Ub12gg69DY/AjW66GA3cYttcAdjWkUXv6Kv0AFb7jRKziwh+pI6HnUP06jzvHn+
lqI2fGjrLfBWuXNg7NpdlVVHpYJRP28oVcMySHkF06y9OwGibgb910FUSVRHbG23ouEyAUPwa8sY
b4A5YsUz/VVG1FWG8nBT+xBDItWoegvwj4gGfb3dPL9UYqlj20ptyb5veEsWU9q/VWLTCw+diL/t
lEn+ToeNd4eItMZb/+vs07sT1wzuGTBoF2K3bKlmE5i0gNKz8dFrqMiXFY4M7HoM6RuKM6Lj9s43
6o8rrQKuT6fPu/dkVaAGgMuZPpsiYLpsYjceCeeGrkfdRKiMivez4paZxU0qTVZjjCe6IAWJ2Xkh
e7uLDtHEUnS9HQljxp77wULCHUMxW1xGS506t913i2nyxq4LfAgnI9Iyy3ri6e4VQeL+CTZ7kr3Y
fZUEEavGusL1Ned0pGOOfQiSCwrkVE1WdNQ3BdHRoigh2N+PSq1kVsmP5BVFLjAKYMGIsUA9uiAY
zLE5o7oTorEkEE7Acz938WmWhBtiBAcoIZCczr9sVEoRqqEUO5QomGDfQj0b4oh1eWHjhSzjRP06
dvVuetbMN4/n+LaIuIZGhn95qnfPZdVplF2vliCZfehrD3gJFyI4EbnyY/XfPpoDs5voilWB1qNM
fAb+QLkvI9P+myIgFKZ5E1FL0selxX7c2fzsRAEzoMpRd+J8PJGaszyUEC5MVBqlBlUjfDsGBAdh
kjoUntbhutd5tkJXog2ILPebcBEbOmiqjRqaQHy7IsrxRyvJcBn4KRp/fHlP57+4m5956EUtwHBG
B9S8DTwRjvhVZt+YblB25f2n7iSh5urdMCAsx1DnWtcWftZhIv3cznZaqTDmY0z7bAcv7HbixdBf
wzEJc7WN5f+sRQ+FSjg5fO6gvwGAR1G2WAa+I3lidwMiIdTao/hHIMOvYGMkbiJCcdujtdiVsloR
bZhCFOQxVfuMdezr26Z0OAC9iPWeZwntMuwDomajfgHp3H1ftVg28r95NIv/bgc3yEc3ckr6zm8q
DmUfXIizEwxGe19K0cbW2IFIEfbORK2Nn/Ad51FBRqj4GKnwz/E3sXq9jiGK2HBJrUDq7HuvcwH5
UjCu2RJYKJx+X15/bSiPeSiwAcpdoZLvqm5VifTKYu620l1hMbwlemjORzDhSH1MKZG4kSMio5pw
Jo3RL8JD+UcRlPI9vcVQFxSGgvblrY/Z2nbEYYJ1s4NxL9E38d7bCmjFUMHNdXcvTn8FnpEjpGVa
OVjU2s6iB4mkLE+C/zIVjnfllVtgJt9/Il3mkSbO2vIYJ20sCwoHotSF9WLYRWrIGbXHY4WPEkX0
XOMtQ4v3pHAnBivoHLQVZgpN8w1/j2LOhHtIStPPNQAesofIEGbwoNLxUKWusH4KtC3S2+5cpFoH
MMHf5Cyvya0+Q29bdTHi5uENOma6XobL/7tklhi6RHAha2Gkat7QNW1qQKixmUcMxtZfsKGA3gDu
bpv9z8onvU0s41TlNSVgb7Q6IsQ21Ev8voIOaUJZUJa42Q5CteO6X8fo1kgZwrcRTZlSd4Cju3Y2
/guIjeHbXnNF9zTg9vu90T9LML2en49tRZQzM7Jp4Rwf/KnoPmgtIs7r2bG+qTxz9uxpzi/D8UwW
9xv3dCtVR8wHBk7e1B2//B/mHOGNaEIbUXewHI9xS05bcM3ohzQ+akHBFARLAJv/fZNsQoMHt9f6
WeSIG7tucegq1zIOGH6gozg8j7HSQl6MEDqp8UpEiSd5+TKfeDZSeksLdSx7n6jqe1SQ956wT084
KkY3stS6aAVmmBSyiG3nqmqE+cPNuEQjuP6Dh/A8AwFuavrFxn1tL6wK/m3sGPg+6YNFIpmcaF4L
jBwfFbO8Frpv07NjSvkD++NYBox4+L+Po8ywFY99JuNruWI5cp4ZFvEx8dhJlMvSjcu/qXj/dBVJ
/g5T/RXnbY5balAs8QxkkNueI7jdQxVSKOCKJCeMopz02zAiSgGt3cDnyyoRd83IhhK0f+kppkZl
YopeNfQUMEyLoxRh9VgZO2Ql4mC2ZZJ3lMHACykt8x0PqtyZC19hE8AUZqRwgylv++2M9RXv8fUY
0CTV+ozTflvFBCcKRog/jIYfIutEHcXlkg+tRkJ2HtUj6pxz5vqU8woKe/CHaDDNxgH52o1cxLi0
+ZBteg+SFiTELP8rJ4etLpsApTGoiuVYHsCKetQPvaKbc36ckJovOp3Xh65YvpgY3sOULZvtXtHb
+DdpOHWcNJeA5rwHuWN8QGA1VEmePUrmurluBsON6WTjwTLy80m6qeBgsq0wQ9uL+WBeWzwccKlv
ROLP9t68/JKMfUqN3wg5C+OnGpaC0DZircTYb0pmyjSun0TSDrUsp0WyhcL7xsKGn7ZxAs/4dAC1
kac2vHi3hXJOo/zwqBZf7tUL8BjUwQy3Ih2o0VjNTt+NaVtG8B+zUxP4fQSqSyS0WHpNxKXe3uYh
6Aqahi4thnm8TFoOllg9LSdbC0tJ71sUkuGajZMWz/gnzt+XPDibwrmxDmB9iZWtnoCB6o9igfxH
YNsZ0T4VPK6eSFB9j8HbdWR+yk5zFTh9Tg55d28bzRqZkDEe16U1LBNE1qeIjkH8hHIEzkDN9oXL
xvjx4pL6K32okJEvJXk31JOlQtR/QTOplCBxw5dtvjcGNNJKexvwtJnwsDMeWAgFNekDC4pKIssm
99meDZzEKsm7ZI8tDlUi0PC1SJJUksrWdmixVD3A3Hu4Jpu/aQ+bc6aBKOWRiXowbXBID/q9nw7W
4ItsLn+msLxuens5fS/4WcZbR8WZnYGnNZj0UBmuYYtnStIuV8gXeUPmhYObfcjQRJgCROPjuoBS
04UQkLWcpS71O+qq43erlfe/r5BhIWBKBX/tSuwXKvVx1IFqkYoI5SIUCj3u12WeaRkbQJP7YojD
99IO35Mk6GLVe+28Qf9afeGetA9Rlh8iQuiN2CyhxnPe/67KujGmh5eEZaFKlvi3PhYbWYgB+gi/
+0YVbYgakBR/N/NGUfy6V4ifzTP9T7lQZvpdtjXP2wsRqAG3ffvBXeBUuP4MIB0BLxbowMgrCQwR
r0yZ2eVsXnIKjOwDbpCpILafqnMrnUPuDsOha050qSATaZzB1AEoHpRZwEr6WFqga3zOcfxAhb+P
FBu4Uxg44oIvZbC50oI7F0ZXw7adcV+dssDtboHoXlRMAYgybXdUctB1YVlea6aKMvJOIZIoJ2Pb
79hUmAJeGIdd6uUYIU+tpO+XshZ2AIfcUWNm8XMpFCBXJAMSNS3GsI+cvJcyu2eU9b0ElCSAeXmA
vRh26wOmVk6jF6PzCRA7WqBgVAhXgdnvinwlMHVCZHSBoLcF0hbzf+tQwd4Yx9PEUh9JQwAza/de
4BDGSxO4s/BZstFBbUnY3BntkZeGioFFpWozmp2HLMBhjB/8EKXkuu74jV8u3apkGKLK69t5C8V5
Y9fdu27ddlNDKli2MgOmxoLTVW4aeZOpaj/Sp6XBRjGqII9ZSVASaluCBTBF3YJOk4fxRpoNrSro
w56mKuBATsoizp8kdg5ySmfc1fcQXQLdcBqrivgz6tlsp2Zjn13fpGAMH/707jNe239LySHVCdS/
QsJyrSdK6v8TPNG/Q88/vVstu+52sSM4SBmHbFIINVlRq9/nuyZDM/XKtElre6UgDkoLkfROl3Zi
lr8SpMHWgxGIITLChi3l9niL8lKcUU88BzPd9tIXyPmObZNVtmq1VKKulLfe7clki29SWXTdTlo2
r1nvHeujLekLHOi6Tu8u6kfE31mPMc1cIpODJnF3oJi4bzf5sM0fQD+RCxUXSADGMfsi/NA9XMfT
QYcssU5sGYYTehNiDTPPszTjTBdQ3ftAqs6+jdWy/zikHCqWhsLCrgLATWzYRgEiHIqZ1RXDaVkH
+Qd1+LcINgsnpqjSw3+OVPjSPtVra2F2CPqHjZFWDC8e7AnpjLizaszC+Q5D+Ybc/i+TalEEvNlu
wkLWm4OdMaOqcyh8vIyyhCE79v7RxnIVbwr3R8pLqMU/ABC63nvcyy1gDGiO/voFVq4z7qr9xudW
v38j7IQraeR/hvs+c0RrilPL8/8VYUdAH9ikuULtPmI3854vUpClrC2jO0ZBWlc+ww80lym88fXw
NbimZerdBosRgkY3q2ROVy0QH92YHr4eiYw7npYyndURGGwC8yb94YzvrYTbxuBh6elrbVDtHkhE
yDgVgFXiAxd6zv+my9fb3P6S9iQm4dfFgqIdo8zpfsY/67E+AFEwoUpQTKIn32FMNHo32eEH57Hv
RJC69VfCl3yXFwEh64xkF6zjnYgPTLIG52bXRNiKTDwVuXIBexnBM8NW+XLahTDjTfRkCpSdYqA2
DvczDpHq9eSEA/mS17zDmEJvG9C09MlVN8myIbrydvFmT4TSa5NprP9qTnVRSU0ZiZKZ5Ep6CPIj
X0w+6VXtU3+WRlqR/Xks5+Dx5ZBF2jAB4zQ50YGV6w49wj/G0wq+YaR3arA2T/dbfq4BW6LkHjsp
lvGxmetIDMaMS3Rtdl+QnZYmxuJ0VaD7ayTot55kXSP9itMOVK9zeKZgxwvUtB2p1ZjuXxlXeoVH
XhIq5zQrX52w9Z0Or9x2z/pv7yoW/au11/JBROWjjKLI7Tcs0VKN0on7GcwtEQi+CKwzast1vYU2
+QiWnenwq5q98hsTCUlCYdvLKI2MTDGSAKzW8Jl32RMRFmnCzbS6c+Qi9TG89VASbCziWPQN2ZNe
GZtZKv39pc/qCsWqzdq0DSab+1q5jeyLlNbPO8Rfo3JIlScZ7NPq4+B7kFIOg+RSrV4dDlL9vLvf
zh0jdycszy8F9yo+nnSHbXnO1j+R7FPomyrbdwSDE2YuxJGitWRRlIAphJjPS2rErkaPRJfskjv4
8EPFSuWzYTNXpL/MqtIYW5vZlUIhXxVuYcPdvShtz3yJ+erVhNJTCPROMeJgEj6mq0zzuHAhiwtu
KeSksXWgfqoBTs3YfoStm+ZFxUdgIMW3EIJwba1YfY6YtOCF7gBoVcUFj667KDjvBFrgct3htRhq
KvGr5o/lv8ph7FL+heqJnS/5pdybUmMh0ld2ahky8D0DhzY9eREO9i4Fq6NVfmwY52fr6ooCFxim
tql+nMT8IT29F4PrymoECFGZEJLejNVcsduvnQW+cjnKvwFtYPtqw7KCyAkud24Cc1t+BlDbr6JU
5nAWk0HZ3VhjuG399VgCOcatOkbeVBNoEpbwaufFvmN0NqsExtlKRaONmPvspyH9X6ZkCz9DuByo
BRBHaJW2bg7U1eSyJmlsy4E3RSM7jpOoOU+JvANtMD/Dxt+uOJ2GpAHb9ZzlVVFTqXx3W9jAx4ii
ozeUYdHjExdaF15OW9wVTCKsfQae3wfP+Dp6QyTjrihaTeVPtkpJg1PPl46IY71Atnan9zSWXsDx
EBwabLFYdE9ydoc7Nu/w3sY2waWto0xm5DOkwtcXARVwcyhnrWulUgoU5ZInOuJaHzwN1pIx9rtK
790ijwd7up7MhsNlU6mGvpYbdvQnari9QedXC6Fp1JihfybQ09EEyTs/GP9zuOIZ7q9hyrGgHhpx
1H8tEwX34XObB3NYuMkyzs3vAOnciclWZ6dxiHo17lsDJO+R0XRKC+vMmhwmAVq2AbwFS+1RThR5
xZp4Zw50KMf0GDn/8ozNHSytwuxDO5c5iT5fuk3I5lqoGZpchHYe+Tal9CIjwZcJbvedRCdbuDAK
a6HrP6S7qJGifXBN2zW1PByL7lPBzT2MI5RsMlZBNmEUd6HjpJ95rpaz7ySQnC5hnrGYWw86bFrj
FhRq32j6EeYI6awMurwLZwMfK2JQopSc/diRC0AZC9l2t8LaCQc0ONx0q3S6Zexm/e+AO5PDilD0
touFWbMrSsb1n95VWhVerb+jUak66WwIlMMUg/m9oP/ySgOym7r98K8p6Si6F+okjUkLSyA3Ytjj
fYXG0wka1wNA3u+LebLmO2TUlmNrubmSsUjkwqshTFIKo1BxW9TpXoennGlOkdJlxA7mELu99a6A
BzLN3T15xb6j1Zb+lpfW+Mt2nXh5huGKEUFej6ezQpDD+uKlNS2Vr9VLgKwr14OQ+oYyc+0BB5k9
CrZwoz0f9/Ss5wMV6pcpcZGNL3p5gKUV4JrhUZ/uEoP73xrgiZAsmz928VZuOsRX+meQ/CqtuS6X
bORztVn4yZX04heXXtxG28chy/ZT0eBd+IlHnf661cMOsYQQ4Vur39kEJfrEY0/D32vUimuWYUcP
sRPEWNwgjxMvEw+pjtHEGhspxPERHQU6T8QsSMQivp3BLOFQ5jiSo+bUuvAcsAAfAd/6zzLu9C76
7Y33Gyvws4fTqUJCvnSbdK2/25kgDOVvHSvqlD8SNeMcgGqZnPFtKTFP8KtmLEqISiXzBNP0wT+h
T3yWcyctNtEw2ajTZlXdiwJKDI+QhqCJGlOtJvk3KnFljbX8YSdwcuMjB55OxLv85ZqdiAq6MLa6
u25yNw/ohNuD4zDfUp6+LnCBzmtmqhfpdzS7lHs9WT6fQ1lclshZukIuSVjpFZvPZ6TfjEMaKWBV
EjuASZUewp1yAz/o22+w4suJYmU45eZK+HTp6SkXnN2oTr1zAhoyqablwJpjBqmxYpWii9Sg+iCP
o3Dvv3DFTUGDl7Dow97OSadojdS2bfGlPrSJ0z9basWMhvYXCzRxXKQ0baLxv1PYfbD7sSkd6oMs
nN4ZjcadJ1acl89rCG56nbmM1bGtw6iABZAdOx73+4z1v0ENNtRdysg4MP7+g5B/+1w+MxSrNNzn
THbPNg8ykJ1xqxVpambwSzn/L8sqMj2A48K39f1rtNpsYNPG/0+iLXKYLiGPgpY6jz39H/gm6JPB
pdv6YuTQsDsZz6sOuFUp5i5HVEpLm0F23j0GD6Dosr00Bcq+Avz+nFUsze3GErZtOyC3kHCgEVzN
E3hOl7RJyA9zW1fOLpoD5UUy+C8qQSBKcA++CW/6X/jy/hk8IO+fHfABWS3BNWcVwWDna93BsvN8
C4EHXVaPotRappwt6OCFlH2KS6JzWTlLHx+BsKqN9ar+hkZckOoI+n5SLKkcPLCAzxyXHzeaT7Ob
GHi0ELUCVKf1B+uZiGyGABp7ioZ4wLHbg3kGEzYRbqYBMfYnqLJlc7qvHRi+QLRYRQvci8HK2ZV3
Iozs//RR2IYJDN+zfM8TEaIAw8unG4C1DVxFj/5vGb5TlErGZu85Gog2pGWNj5wzKkis7VdlmdB3
f3IDM/O1TKPO2AwSj9Rua6KQJaRW0n8W70AuxkJJNLZWdHgmjxO8sSZ/sR2tS74lRV/dKG1azMs6
ev4y0pqWluSivEiFltK2DyIubgxunHJdm9VCj4D2KN2BI4fPEn/sCOdmtTOG10nN5Lefy7eVBiEP
WMv4ie0rSoL0T/9IboGxwjjR//qjuz0RPaGvXLKdnTCURDLM/raCOWZRrsE78hHHnXfYP5uRKvKy
Wtp4jum5ZVgmnLcJlj3PEXlpswAq6tIDwZypdchkB9RQkv2ygPVRBxyx0oD46gyTRDTdqRrMcY41
dR5Yl/+y3Y4G4P8B/HntLgUsqK9//nVI4Ojx+mEGqzx1ui1dPYNRSgfsWm/RnI9bFawJOYgTqz2V
+g/TuSKXA5KjhqNdKnsAKgDgjo73xazmS73VnclmMY0gs/+Wp2zy0OjQTnSH9RNWQf6g/6OjPo+G
EfaEHlKh6OuO59SIemUoK2aBQkjnOne0Ac9jOIMcb5T4X+84+riJfKUx7PVOjhYHYPdQ4bOWT+2e
rJNRaYjSn7svmldy/su+E1B5Mqz55r87XKwHE62fZw92LyX/e0vWlGnmx/l54Q9xNV48TU8sbduo
T9JkghpJ73uKoqSWp2hbu3Z4LVH1DnNVySWU81Q+IJF4URj9rDzmWaM2y4QGbSen0p0Vfc9TfCeP
VuqBpCeoP1w++t2HVDRnvJ2VqlPeBD7XWkpC5eyeG+Af135mLAR6914l7v/5OB3wnwvNoeY+CaPO
DA1Sgu2JGqz8HC9+Rc53VdZNTU43NpM5eBT++Anz3ljTjtdqcwhOBqo5UuTueI6VT9gT5YaRV+Im
7F66wT2Ws+ch/5GlCqZDwM0ZiPA+h1JNeUkuDVv0RkeSC1/bB6OIO8o9/Gxj18JL8rP/ImVt0y6z
EdeIaeCiKU/Kv2UFwTc7VIbJswJJW3O+e+XZXkY/xzY6+45clvu0Z1domCCCgFPpZD0YHcCVJhEh
t1CC1K6PzUEYas1Ak5kFD6k++o0nAaMc1Ib6Nrqln+ooG0z0NgEFlbPtsIe2ZKQ7SBmvUtkK9fuw
KUQtafhBADO/SR+aXmuqxfsV4jQvTgNIc/8PUrYqT0KCcMsoUeQkPawJnk1Jn73NtMhQTnW/dGsL
wKq7ArPjOKNap47PUhhhX9d4yfgb5+teNjoUjWF/t/H61eyNIoFe2nsTevuqgrUS8Q56ZXbLagZR
2rojixLUAFrk3WbiDC8X1neKXZaD9PGQFG/Ds3/i5YIq2s9OAs48fcmzHj/ziABDIRqr6I7yfXOp
gVuHBL+uF7U9uykZLjodBF/yCDeCzPvkjNVZR2XD7WZicumWKDDWBL5Arc/72BYu+AqXoiTDLuKx
Ga91/lIVrA2uifyMTe/bf+PqCDuLYwOS8qMu5gaShL7c3yyHk5ylepzj9a+aNaJtbhQ1qIlIjo4+
SaYbII9Yc54Xj3Lch9GrMNpggrjNpxpHiAIxyqej+FM9WLWk4yICzxWqXJBh4DOS9qTCzlQkF98E
Ge1Ax9o9BBajL3gvRrdBjLg/iM4oWmnN1PcHd8VjJPbuOeevQ6rA4zoVUALLRCLQTDsmiSL4qjOV
GzxnXTpqMOlMumwa2xFiCu8+FIaeUWHhCkMisTJXx/80AvetC7qNZrVoKdU0X05vvWadkd7IHPSq
7+dQK7QqkyY6Vbl2lmm+EAQfuDrBy1viV1at5Hyb9X0Ilmy7zwJuIjgyeddsAveFjf0VeP4Q1krt
DGn3QMgjCGy7NLvM7HpGMjMXeB2tQVZDgewcA0EPhd6AigskJzRt6i2s9Suh75hpjgg133Ns0LIP
ku4jxFE6YIjp13YQIdFG6rRM/r0RURksobIEl/tZl6jEAGbql/oclPlwsjCwKTSsJ5ZOFeaqESDE
lOMvA3cdgV9rDJgOgK98G3ab7WDytdbC84xO+wON8lOnXxPF3AbaBTjHEJAHtP+g/SsiLkoO3ZbO
MnRijUrt6v6PTsZ0Cj9NezI1UmpInNmv0bMbcTx0cttVldhzgVFt0kIU0M3wsCTzZPFHqRkhbokF
kzhonaHUJAFUPfC6lkLHuNF+PUMUIcjznitL3qzhxDhtL9N0fOBV+XP8wfvgs+eRdGoyWGAgM7Og
E305v34R3rg+SRtjyn9eSeh+6HiygkTczFOwODOhi6E7RYk9ZBPIA+sarHw8tanhN3Gs/H4XFBDr
8z6kGCXqBb9w/KM0a8FRUPFuHJgg7vyN7YIZ/0KEulVgiIKq1yOD+9Z8NP3LW8l1NgSeuReB5sUt
gW9EAIkmzjJf2gAqTynO2shNoW353jIqg1QrYzDp/8Lc/bh1oXcOgmykRi5sHj9gQJ4PDiepXhOk
ZdGG5xhqiMl77s5zrhJ74+3GVk9FtKKR+dB+g0k1Ty4OKlP6KSieW1x5Zzo80mK+RcdVK+34pDiW
MIR9QUhLrHZvSugDGdCcvhFQYJqUINQB8atVz1/vtbI+n5SUxYS0xJoUoUkF8JVNjPYQSj8w574I
pcK1IvMZCvIxuzk32CZQYilXSodmY17XeUdexERSlinvduLXlG5AYB8zXqQIXkvaX7GJpyXxObEg
9nvXvwF0BaZg7Yhz/BGv8dBZ6qb+QtLWz446tZbUwg7PHIGpstXPt+EPXuOLeeQj02NuWuttsCZC
vabbNC8iG3ST0XjqJxAElbQyKmGgDXw6ktmQnnDSKcemzNJwh5JS8v2vkvW3WrDak2drwxV26Wa2
y2tRLuV8TjbC4QZzZk1U55gyOUrdMbGrTHo317PpxwqFV6wY+qam/lb5EwXxNUkHkg3A/10wDHnn
5EG6kLEx2W2alCpYOnA9SSQllkJ17oqCe1Q/2ulc0ejk/o1hsrlsC8dLRr9yFuQhR16wYyxJ3UTU
1usqPfJSsdOjWkJC8mmdMrKenDxxY06nyORLtVm/LXrZCH21/w8CW4RpaZ1N+iKnmG5QsDz6kvn9
xtDAQzgLtCzIhB2LjI9WUDeLkFEjslY09liWKHJ7M9ULZofPNUOkcxFp3ZnOn7DuETl/AWvqu/LE
KDqOaBClM0XFbnPDYGSO/10eIUHmbGjuRHcOZsJhDnbkrs4lHQOrenumMr9kNEDNONXy4/r+m3YS
qVhLoZmtY4AqOtJ17OiwBc8Dury08Ovk4QXX/hS+qLsNkj0l4HBc4IxzB6kRJ3f+lx+b0YMFyHTd
t/OW267rKD59VfZxIlR7sPMj4dJPQhmxzPvmVgNsZJuSyl13VcaemUlVzIZmRuSPb8gLvEvHkWXG
cNhCZ2fIocqu5jXZAUc2pHPnAU87Qtan3bEVInQgnhlx7wXast28xaaDvnUAisPBnwxBg3XLbbih
4B55R0EfjDCDB6TuqE1bCsPofogiFoYOle7YS7eirVnkrJ1Y3dVgWbr2kKnH15k3q0wbqQzbG6Uc
Vi6itVeidaXjVJ21Ut0hVyDex9llWyB/HGDRYeBXVkkMbqwcNu9yWqJVdK5acCeWZ+gcBG7yKxoH
6fvtvbXiUi+uklj9F3+ykwY0ntXecg3Dyzk8aLIkAFVYL+s5Xmw0wLRFVDiLlfASNvWAPMc0Mv/n
OHHL1LMfgg/h6aDZY7CyQE+i6bK3cl60nIPhM/imnXxfR/1RKXzykbsfl5wheIR+ynZvQLaiezJd
cEwXpktAxi/EKBgpWRcjsa2ykTVfSWQaytd3lWzlhBRR/wks1XKG0Ckld3L1No/DNfN8U2yUTOgS
T1HNygHpKZL4SZmCo7K7Nw7SMQ8nYOekdXp+p850vRQAYQQfGybiI627MYssG5S6DFIUHUH1z2/e
w8gQSo38DS33Ahp6skBCKZz00F0UzIf8Ip1i7soBSVno2Qgn5xsREL0htOTm4RNqiyCDsrO/sRWP
vk9bgTALidLq/5I19DRGct2FnJhBHBJCj5ylmfifDuV9AdrOcDISM5/Q5LZUxmH5aYo3PXdsgW9A
TQN1/2C5EtB6iM7AEPMoUCVOvRBb9JmqB4MBv1fHWYZc/FG1kOt+UxOSwJJsC0TfuypiN6JhtiQ5
6HWd9Y7nlpIvo8Thy3cDvAC0qXOsLnEc4TZLdft7hZaQWBpeq+U1KHLbNY5IPVYyfS3M84lRDHq4
mewTSC8Wv/pdAJ79jlwAWQEeUzFZidivnZfhVCEDXp4Pnil1d3PHXs796f6JgNBUzgMIunISPFAL
9JlM6WRk2mqawI2roHMvWLN0VLtCAD1wkqJuyQaUMhZ3KAAynlp2uNSVm1Re0JN66Tph6yhVG3TP
3OPSzDn8lG98fD+1DtaITdo2wxFc+0jq7ztmzsH8YkDwBkmps3IYV0hrkCk/55o46Cec+rmPmRO6
7Ybsh4Ktc9lWCbiyJull/yQP7dza+NTXusBkjdo6QtgbqrxZHflX5k4uwMxiywlfthwmfEn54dJI
3Dzyrosk3D15chWTi8SBF+guCIkhwS46TD6YB4kFX31dGKkjQ+Vyl/g8fV73hDx2umY0WPHqPehT
izf56oH1v6vH/QV995YbTJ6r2M5aeM2PI6vy1yfhllOaMBU2bHvNLZQQP0GAcuj1yvDwCaHxrwQV
VWquRuNxqPuLwWgn3umQUf3fpc8GEkZyA3VxjcHIlghehMtf2W53/SzDI7MpYl30WkRO0FH13Wgt
VdTT1LYHtwPnWY8vhouEn6QG7fdV1WonQtY+KbKg+mP3HxvDAFJF2zN73+gNZ/gBhBPMns4vRKjt
UIjo6tQPg3D8GBTa/jv3QrUUcgCMIVowIEW8XmHvHCcQH1sDAqQ+h0qTzx767lAOXJWe4PMpU+j2
5JVkCglPWo/2pRhL8xfMtesoKL7eIIorzmggNN1RDrTVUMg4Udfu04KYME+Hm/eXom7yL8txnklL
HD3w1va4yTwTjEljuCH5AiqPNbxlZnuo8p73cj0VLRSfXAyxuD1IrYkHpQ+vikiRurHjuPah1Ec/
2FQf+3tthv4SiYBHg22l6WkAo23PIoMXMJl8sFx9rwQ5dvZzSJs3K89oOtkydyB2Rt8wwVSz7cmr
E7VwyvVsLJc/wqPWE4LE/wsLi8fqSDWNpr8JUXfa0Do6ionmDExTN/JLxjowphc8kY3X2M+5/DMx
4yuLGY4F2nNcMRZ8GIsFCStb7X7OVN9YGNsWgJnnkctqVODWPd06toAFffT9DSd1HY09uLNPrkCz
Ed86cUTy2w4WyOE9lT/A6OvvSDU2c4tdiWejuKylnE8JxEOZlxIz4eQ5puMc9XIflql5du33ESeb
2PUrcMRn131kgfzEXZvu7Nj8LcOyU2RQAF7YwYys6HjEUt7nPufzug+6Nf4jbJvMqkoWYNt0b2Pq
d72HftcA31fAymvmC9P4hvp8GLsFElgxOEbmKH2mQ2SxxaGtLp6yeUuWlonXMH/Zkxin2pg4XvVK
H5jwbgKybXoT/CSP5e1s2e3nIiiuvaj4rW0Pat7INFAcV+Uo4uqpFrmyHfUo/yzyqQxxy8x2lb/t
gwm6tgISzjhCRjC50p6xb7VFd8F/AGj3t3Km8OA1LyAgRN09aq6rU3Yx6I8F05hsuC50C4oWD46b
FEV8hSD8kJHkPMATXbIsSJW80DPAAp0iS1E//cnBg1zklx1NHMhxvrGqD6+ZkZWrh2+ynr0Ozjjk
gIQMVjTDJxPgZIkgmFr1v8owHhoZwIWaQOjezhzO4E+vku+JGCLlZKRb7dCGCeYTSt5rG/dJYrwm
GHKuGvJgKXTi2APVIVff+n5tCd+hzQPRzJcKHd88bwu4eS0AFtDBLy3miaomDWQhWcb4mtRXSbu2
Gb3riUzw4X/R6hCNdHTBef7jHPvExAPg7G84T/asRLnLiWPCeCcxAffPrxOglA2nRd2E+n8LJR0w
dBYZ6FIOybFIzSg1pu93Qmcy0TvnwV+ww0WRXu7v8iF8Bu22F6YKA1s22dGltu+65Jq1BHAG6SnQ
sp8qNwUKraR1oA09pCX0lZKH6i2pi9C3OZuClEC76SsNXINXSHE7jUD6kjBFoLwnFcAGO9wLeKR4
cQSQQdtm8tjm7qtVHqC8kQr7ydTxLXlb3oGfpj65igeDEF+jHXWpC5NIKLmopTSwECJc6Ki6AtTi
ozRloGsx/ECSK6rZXEoKuORQH8EmEvt9ghXpBTSySYTidv6iTx4Ect4MP5KfVfm1rucTu63A4RPQ
xodQvTZ/NbG9oOoPJoYO6ZOOxiBx8/K8+7UyEwUt7hquGXDu8Q3LaaQjKUmQiK2VWMCc/unXKgdC
Wqj1r/TlJ894ztJtzkOcVa4KjgPIllKMTI1nHe/H7p/c8UjWTw9bf2/L6qqbmaFVIgljZ7ZyBQMf
XCNocAfIpBFkK1bQu3r9pX9RLWkfEY7M4pYnoA9aRX32ALiyho4Eise62Vc9FL9ylhrDfkO1oA7o
/l52GdVp6uENDoIKcIT3oUg00VTguTqyhv1TAr2pSOEaS0hXTeGPoO6tHBGcu1rK5yZ+lBNumcMs
O8ruq58a9AfHpZAQHWOPbBbfGRDF9cLrJpCfhJNURktVi/MRub3VZMuLAL/iUs5O4AL7txBgmbK0
wtzcF6sangGMcgkGnl+QoJJKCuu7vkvrO8DeSG6zofTngfPY3oPrsteJxY0EgWt15RED03Frafw0
wM/gO4IkZiDsWGEqwlFdAmJaFAUbibOCNDHJW6wRoKRwmI+UXUEJb4epRjwRQ8TgZIMzIgwhJvbu
JL7KldOVFi888ptMphCX6NCzzTEvv/VAmW77doyFg3524JIMRV5TBAdouKaFhQW17oeDwVX8SwFK
OxFJq7OPECgrqOXvHxPdUKiZpAliYQkxFHZ28Gjf9n2eyG8KI7kwEMas6aJCHY5O0V64YggqpesG
+PgvZsevLxgIOGeQqEySPUEbY/v+dS+0ebopbVgpcSiDpBy/nWMfO1LxlN5ZCt2vuZuMYZ9b+CsA
OWwyb/HqQAoIamOV38x1RCmxFGHm4lLjOyGxREr0qQVvGRXVd0ZdguGQrFzAdmE3OmnvJ7Re4+oz
O5BsMl/7981wbzkBUfuSNEgMUdXWzqrhKPhHjTB5kiOi35lO6jkhY553KScR6uwdc8QGcTQuAs+R
6pTf4KY0dqn1Zywl+UI1OnxmKjEdKVqLKaYsWdyMTkUZMoceDyQJeens4QS6kGndNfA3iRRlemqQ
tTyfnJXvBiZdWu1+lhbdFvKI4kjHQQJNE+6Ehomw1c091EMMsDLQj6NeRdx39ZixYVNj9cAGt1bj
ZiJI9OSMnFMeWqX/Hc1xRs0AwYRKIxPHOG9ABXShU4DHECxG6UKg9M8Z6Jd01xLJo6wCOeJj6tZn
9o1Jhx7YvfuW8lzKIhffCY1Wt8oo5fr2RcEzt5m9ne1OdI0nG6QMjxJpWxf2TzJlsMHpO8kUVDG2
gP22UFNnJT7xbpyms+OXj6OwyglZPu102niEls1wEcVWZvf42XQ8mlbPZhGfrET46von+sWisfse
D8qoNkpW/xkl9jz1V7o8xZLdCUiX9MHhFE56KAOaCM253ehKrGMlFdvoLTV6wKOSjYKUJpzPLWVP
N2PyI4il3+orou74DNcea8XjEBReazZKwGSvpMFPyGZNHr94EEoPQgksbkrQHvBrYUoaV8AP9aVD
6XNwfK6mBU3ttuze+urOeeVRaJmmI0+mKkEjOy/B7c3kJOABCL33NLOguK+RZcyZH23x8MReZzQK
06in1QCmuzt/LGm6Y1Wai+NLVN9CreSLpttNvUueatqdteydDJ5pK70Oee5op66s2pWO8YYwnEMQ
jKVaZLwCdKcpwIHw8bz0yRZ2TF3GGaHNTEAIhg1uQxYCwf6qtTE4jOluKRh9S80KslBNXR9XGegb
aUx1m1Jn5nx9yDC3TBxvdxisUTX4jw7Ip2UmQDNECCW5oW3eyyn8exoRdsWeutWsJ3fOqKUcSxIA
6Lc3zMB6jujOSUBSQS6Z0IE0PmqFpS9Wq/GrfvB/mba0NDZbrKAJlIq/J/O1yMlyLF8JsQXrjGLM
1K/+avi9VKN14e7DqixoV1H5PUFspnPW/hNQMSlVK7MHvonpb0yIik3OVjCpHQ+vyM5kyl/RV9E3
YMDRxAvCApUhHpueYyfuOANfXH0jDFLJGpAHMbJV7Ag3D8owvETIgECBZEUESsXSSozcRw5iTb6K
Cy6uGna8Gx1uYWWoRftPrCeLFCkUywdZI0Kw5KuWVNnR+aMlNyy/aYu7OqXzuvLbGNrhZLPz09YY
KRLRHE8LSCqBSRxyPBxcF+gcK72Gf0D71vYGd0QgzQoon5RJbE5lXW3DaBqGQLmsAyI/risd/MVQ
yxIbfth9A5zl6e98zfIDXuQ6CJ4/n798g91canYr6Jz346nUt8I44UVl0MqLcFVlqtxbgCilmGfh
QAsVaG/HG5S+aiV8yBmTXXjvGJS3erYyXvDrMMzLez4r/rQxMi92in+CZzNHrqCvAnmdD3gFoTOZ
tFafHvTVYiDrwwc7BbSpE9TqteumMGvQeChtcQfdOs2FCGNoS+7z8OJjkukGyzWwP200vYO/pAsO
ynfd2emJvizFS7nkdph1dqQpIftwDtTMyy9MJXx89LBQUibsnkaCwblbJ1scSZM69MysRT5ge59t
TIjPCxfqt5qEZZ2X1hn9fVtM1iPHoTFL/cH/GNcghBJOkv2vgVyQlIg2MqqNsnw5U957OHvlWfc1
lT1c3q5dr7ylDkTAS0oPtU7xSsU54NTuSl6EButeb6MzItOigv3Fcho1NMkJyGxn9xjmsLuL12gs
1UX6TTZJK7i1iFDl0hmD3Q7BZOf3dwHA7soFGQxHYZ9EtoCVxctsSoqTb4uyvc6DvN7LT3lUb8Nz
GdI5d+TbLSUUroAKX7BiV8fChr2CETDd3CASRanhns1j+tWloBoi0Q/Yw7kioZF/AQvE8oJd9Onk
QLIFet+W38tKuo9a/XaRxoStX3o/anxvJTrjkzypYBwR7/OFk7qitW7VOvgO3UQvppScajKvnAZt
1IbwfFOKn3U3Yfn0WsrkRSV+CrpmFnm+hJI6gmwa7P4HkRwMM2hhkD9g5zish3rOImc7fw9q9Zf+
ekKVDUGoOfrMfJRKE5zyLKu1JWSoMPQEUXbiu98sR8xvbqrlc4TaPPB1Z8Kky4ddUkv4bgEBoUm0
fRo4SSNNC9P05/J3nQtpzHadHtAEuHYRQRDqsj/TULEz/zciJGMbh9IRibva3D2H0cYzWGFmv73D
VIiyIiAp8nVLARiZRfzLfQa+WIhf6hKH0Hv6pimxAiDy/R7I7YAUp/OwEtL1sBqSg7OhcRnHgA49
7i+budcDhTf7Ks48B9ihJiqWVjlbKCEbxBPMzG20p9Nn+elHuNZH1/R4s5/DZl+62rvUeQi2SPUY
cuznvPQsy/nKkaLpx+ZlK0vAViNAUlx896M5a+e0yK4m39cUpwQrml3LJDUlVYCvD89D7ktMINMO
IKCPQxNAaFpQP76I1gx6fwvXrzKZychhwBijPsyqmc+fzqOKoheXTmOaZW+SKbYhUdZPZ3YtIGC6
53p3GzPrPSTA+p8Da+OYiLk9MxFfb0KbOn8zYpQrCHz1TCdTGBFJAv599xPiIoJERbl/seucL0Sl
pkf4N9IjNN+atUYx558/7zZj9k+N9Z+IYnXTlYaaxOmeulC2g1QdckB6p0R8rZfNvCSCjJo+TpZP
kCiOC5UrcyM/kM9/8gwaTYi2k+VWIQLsx9WwXYpisgXSSctPU7ncNeDal/zpboUtNFX8tuWZ0P3C
TzLv1Vm/lsHEPPTLX6QHyZ7a2UFfjuAkCDqeIkQr7+OADQPrgQrr2RFcD8hG/Cn1NB+ngznnQb7I
Naucp4R3sKEYmwo0aCJ1W+7fcNMco9oi3ulMAjNtxCAoXZitQsn7xeDIfRM31YILgEVwBlRc+RO0
8Gey4RoYya061yQ1BfsWhOO+T9VZhnQJkV/Dye9qITHHEthdXtSzt9hcLMT1HEYueJnIfwxyQPE+
nmKkfvZNw4gW0pS3VZvnr+eglXKbl4ilQo+9+Qbhh8t/+KxZ8m5fTHNkKrADGYvBWlAMbBefxmTC
Qy1At7jLxt0LMhHIno5OMHGSwzJdNMVsKKv1OmjgIW+YKpjtA6+990FO7nI/MgvaiwmlPBhKhp8z
QMg9XAIS3UYRk1EmBNSCeyAZe9FD2ut4sKIX4Tr5pFrgVoK22hxnznnRHOyr5I8w5pikEmy+mJyz
mXpjioms8Nx5nLq42QZWPP2VJy75u8vtOFESGRGU7JufPxershlOJ9wTW3wCsSlIIGeNMHyTK8Lf
cJJYFmbUyQFTzSGf7ks9adTOz8V+OZCtRuSZ5rhDc3aVyFPAMAwnQN8R4LZZpl4JHBbSKx5ECdo3
/fjltQuMIyTP2jDLqrLfu2146ig2hec9JioSqemG9rbKzQhNcM4apg1vIhHvwA8B1fed4pZL4IpJ
hlxesFOdTE3zO52LC5r6OfDubtndUrO9t9qmfqfZNDU3YZY3n8xYCU5nPdxNWt09qx8n4Koj/9TM
YyU2k0n9who65NehDykZVvYdNJKcfztQmTB1TbNJqFncbGeJAwdCJZccKXKwzfSCFpXX91Wq4B6l
8Dg5svQnEJ7DNcP0LOg+/LaobVCmuxC46L0OgsCCxsqLORMixeIIYxmboYK/OlBi2xHK1EPgPk7L
Dv9NzcTnjwzezbPbO7oBMUnSvwcBwVPilKw+kqq3wQEJSCcus3aS/fMLPAvi4+qQlryZFUOH+oFR
iQTzoZK5Tz/5IJALTz3EAQuVu5mtSerWRSd13t5eGBXM3ptOca9tVUYmEkZ5ViDaJFEwc84B1QEe
3fl0VgmdZIxFhI7re8Mc3Gz0HBhyF/VnWh9FTJJ4fHJXJt4L1KihgdBwsnR806CYXetlnUlM1Qbp
HpX6w6QnsXLnBoUws2x1cG285zJm12imSKJNkzb/AyxuUDierlmILlDZWhhCEAM1gGafqTKWed3q
+L7hkq6MW6I69rqCvUAxXpd6SXusUG31uZHyY4GBLXnwfEp+zwHjejbWNqtZKTG7MEJXdp6eBiyD
3L64Vav1dd8mKd9IGI73rTP82P+44IcFkeQAyOGNu600pRMt4fIkyCr+Cgfj1d6BxIQH8UygXtBp
/GbwNQdIcXFUROHYScs8cul0rNwQDxtIgjmO6sAaTuQhqP3FDye24uJwWS4El7VNAmND9ZbI3eFk
5qzM4/kZr/WKGg7Pfnunr4i6Cx+R+tz6awodWk8RgYzDBJMXtfF1OovIe/XZN7ncWPZwBSRYf0uU
7MsUw2WhTfjKzIgl915Zx+7LVJ0wKgsF3eO3LiUEyV+qJe4gazg6vN4f0EhMXx5Xcm9FrWkgEjfb
wvZShp7xg3d+c8sszl21Un1OeXgjjItdlcqoCWTE9Z8Y5vkMUpj570r1mN0VmX58p4abVq+D5ijN
tDfyjG39HPMKGbpfX0AAOmVpQNFRRM2p1f8WaDPG+/I1rWOfv6bYLyfc2VmQutHmdbf4vtbpeBtY
OATdcAR9Xm/HE77x3EE2UG+8v++wCyLOs4BVeHLWbivQ25/8SjpGVtZ2xLagUTfq6gsO9/6YfZgP
JwGa+tZStXkUaQNIS5T3rB94mMcxScftIm9MoRK3tG5Nb2svHcDp0/RE2dsaycgfXsgH+bujenhN
D19qOjbA3PJMiQ40hgcHkMLLMVeuebnQH0no9n8kKgQa6IAlaeiW1MXBXKbunvjBNgD7EfJwHtaQ
OgO1/yP8cPIpI/DGpBaO44CyowCfIqTBML9vxRSAYhPIjylTEqw8r74xPnvdcuiAAPEc03MdVYmz
PbPZK9CaqwUwbJJrT+8o9j7o1a0hSdKtGcm4PJPsFM/hPveCXEvcaXu3tlJtw0kKkIyfd/8k7wsz
HCx/M3WOp1XSaJzTZhlTe4n2W2WclxehGs7I+sGbAPfxgqi/4MNaSitmAiAtDzSpdSvqWUejwhnL
uzyn8c2hBi+WK12oVcZ9BtoTpOOjX7DqMO5yZnobGeP6dWAcMLQKt7QmD980oW4aAcIwakX1lnjM
vpqjtT40xb214E1LjJO8VQKs/VRBz+B01I6w09nXKexj4v9s30OvX13S7ZChas53v1M9mGrnhmz+
q4KaKwJcH82GeDimCao0UfUVbhaXQLJYsXKmnwM0suV80lcpeYo32qz521pPn3GAvUaU5vDJKAfJ
684Eaxi4b4Lm7a5SF2rHE4FV+W5T508OGtS4B8h7SzyNCyjcC9vZCU9tgfx1D5+m164NXXxgwXeB
SFkvLxP4ECqnQu55NwmeLpiY0n9cTrh6szP4K9wsURzrOfK2IpfC0D8/zfZMrhSIWTl0B8buZKIJ
+DtNmLdI/4m9ybT/KL8/YhpCyV0Z5UfIo+/0yqQtVmGhmI3h6sdVKKUmdQh/1+ObDG26YA2ouWy+
SSV8B4S1T/7VY9KkNycNgupJNgjZtxaV5OGHuKGPY8Y5aAR2R7Jgxn17+ZU8rqh5R3BGJFtpWI/F
P+EPrdbM47Whul4yWkVzLzbKUO1z2w6j/+wRoq65WmtTKJm2JPjqGhWyUrCHmeOsoW39JnGrw4uy
QDlZOZYgss5D+3CUdpd7kNG15k+fksHDWiL+GhSBXTncgUV+O+QtWclXPZpSLMq2yUGZu0MYfpLo
wiwfx18WqWgPQtT5DMGEu4DWSa2JfXCookq3VpfQw6aq7fN2Q6dw3F3h0OXRF+gREHGbAKEwim73
OCelm3ZtGr0uBTuQXoIdQFDxdPnVT/doiYZJ20e2OBPGZj0ZuAlUkNA63G6yNHFC7Qww2HFfk4RZ
l1EUxcgbQpoVZG4OZZLluvG0gcRHrwNR1NtdUqIIRP97jyO9sVNk6q4FqdWjNMQ/qSDJSAJmiDKL
q373XcrXUdk2pOeXZX2gvM7woT081MNNm1mSCg8DrJLPDKdWAtP0kQSany+OnGzDXFd0yoxQOTHc
kzQ2/2/5PfIe9VgS6O6ET+//C3WKHgPRKxzzsXqpjAK6F/FPbJ2Ybhker6yw8jz6cM9B/SnNQ27C
neEvIooSij8ifDXaGSYpZ7Lu+exPLvR6MmXBumALCtiPb3OvMKpdG2w6U4EreBPHNvxzAVAOJZl9
CYE83jPL/5PDUTtc5rZmaZI8zux8Y6Oip0j7lBSN0n3EQGhakQtnJg6fYDWEpvjVUsBf5zbS0/gg
Epkx5msDdRc6ykPIOBpJn3gnjvoDdz0JbptVdFuhyYlnXvkgQuYhK61LElEi0G3kYS5osOtnZsTv
0458OG1VIm1NPJ4pYbnyskjgp9UmIXz+cL92/X1si9beZl6JRZEGe1VLtzDkaqojWSC/tQ5YKdh7
W4helzdvuh/mJUfOBHuT204usTmz4rh3YNUH7jDzhSfVp0uVGsATp62IMfV/A2ooAh/F/lsoKEGK
4EriovGRXw7FJW0BC0HcRwWshx3TYzszVf3WktD2E5mhh3tRf+B4SXAB4RTP0uY1qne/r6iB3Eps
N88CMF0ZXDIR0U+1MYLwMPYzsJw1oYTVmuCCTntgaZ0Ohi1PPQ1d0IIMSMPPBniISQwjn41RvNIq
hACXEZUMCRp/PY0v25R8z2j/dFCrey2EPbzjV2I0JMobM4C+EoKCcD5+rKV5PMOthHisyY1oJLfv
Gqw0PhezKKSnNwsl0FHECYfHMF0oOCDgrMyKURyLcnp0Eec5qD2QNgdVvxGoPmCoQbz3zr2qHSvU
0s2vgQIJbb1vGnnuR1hywKfts8kglZQVXEXppnwjdE0HCW3cbgNCvNGTijGV5yC2ahoviGYbc4S3
XtwdUxYH//W3/qMe40kFmbyIwRE9hvm5kpoFZPR0IiruaVXLsT4b21y5YkaQoQebFNnjmY5Sc/Rd
r8zNu4BGg7cFTuQYOtwm8/VyI4kfoZKNBrnmMSU3CUzspSeFVSvfu1jM/cJt1snE3yXYEfA/+grz
//W7gdNZcBHvXIY1/qtKOy0/L8uu6zrybx9Vky4MoVzEfqqnNZHiKP0qlHX0oVv+IgWi/SFqVNrO
OW4ptGimE2o4zm8UEd9zlSJ2AQtpJ5Vmr7bXiKDcFFWql+3rC7IXrXrmfspkCd86CpfUYkWSK9Tn
K/FNn8iEeOtWgli8LOdbfnr47qgOBvHUw2FanriNMW2vEIKJi3jaf3d5YdyuCvbpS/xw7qr8t7Ic
pzUi1fvDWm0mtUUChr5DNolNLwB2Wu8Tm7lQMruTh/UkHVzzHAyLA+xb7L9uuY5BJh862A28BA0I
50pmXIPNFa7K/cR8SABbGwwfpJvfF+J0cYvkdyqQ4R0Kg4BSIouJc2pYcrNFMrs72BAaB3iLeFtd
yX2y5PttSjVHFHDOto7MBoJ/t6ffKC62+/0GzrstbMxycHaVexHlwtgmsAYrzyZ6ZXrO8r1VhKjG
5u1zRpSipQvrnclNFp+4jMuki6SKwwVJtkKmCiMV1vaDt4qHY1Y5ETQ+2xZaiXfhU8RKmbmB4SVd
bOPDNt/DV4xcU2jx7RveBvDmTgwiJqG1uu91yT27cSWnear0xaKe4AY7hB+2yuZjzMwxamy5d0+1
IgsxP+BK5pIaztx/5Rd4wMAUzV0pII3Ua2TCxJdVijwCxV8NbrwuUgQsJPQNXP+N/WAbzXkURylV
5Iikpf18ianqbDX8b/ITBYM53o2I76EpEub2A/7gsnvx/mCpzru74o0mNac3wV8OrqM/mL7nRo1k
gVy7QwoEZ5AtnzF3LwvW5w+8kszDQD8rMCEoOHVJgB2xpC0wZfUkYAU9+K/gps35gHAJtoQJS7wK
lmirW9XworimS0NfwZrM6sVhxyqDR5zxKlaApNw+Uwpmg4wl7aZgsVWirAIulCtGoYMUpJYC/rxt
sDBs+t7g6ToJN/qd01coOukt4RVy2bgjP0Dsh7misZUMd9869rBPMhTHXLJsRL9h4bOVEvFyTy0C
mCgJcF7U/wadP5lImqtDuq9NjunZCp9JsifXpoCdgdDvdpiy47Z2Q8PYOYfbTfJaiDk72Y07PyAe
ymMTmQFrw9OLL9z/2uXODTVcYQyN8YuHFnM1yJIUIk6fHY4tVwIrg+rFl+q4CzWTrmDnNcbu1fNQ
dXPswv5fAthj5Ck+WswLT3dKbBW8JCc6yDwmA82yDSQQNaMvi6jViqjXBSwswl1j3OWHPAnjAZ81
UVAbI3zT+qIGULhLs0txP33l2Y8pvaxZNrvoag38MNYBsDcKL0CP+CHAJYmh5js2Zn+mPxtEhUFV
sQOVeb/LIP/kRQuy7Yf4HGxCOPk99mKi+/jv0xyB0BJObg2tJ+xHV4qqVWHvB0CLDBYG/BSXgTcm
AJgq+WxDN7SU91et2gY9Z2B3NpIWVMZnAGZ6+qdyVm8RAbFRKFrX2sCdxyPsVcZSxKqUturHxNrT
HOuIPloBfnatMRPaEJIe6f8wWApdW5ofogNSCMcKjwOC0wuwH1Ra+Z6ojcrG8+dCAH4llcGZiZj2
YtqhTzk1kbL7zNErOnu65HazbC+88qGx+ZlrajmSU33l4tL5+2eo/13OTQ1Kv79ZOjANNYkgjlel
EziE4SX54sRV8FZkW8UzY7ZXYmPAvIPnyqr954lSVtXqL9vZnbIMsNZJ6NyBPES0co7RKAAW/w0k
09Y8s24Enlm/26ZGCyCE5KihMJet5LZ8i6fIlo00HbC+52p+aGmeLgsdmoqSpAYmSPJvjhXXkuyH
fO/8hD3NiNTT0oshfMjDYdE86ApB7ZAMbxgLR5DDjeW+Oa9quXVkH7uo9ly70U2miC/OQ9/EoX9m
ze4TQt7CA1Pf9A9u07bVZwNSu4ruIFWXl0QaQbEhixbS8zKGbMePNzXCQFlmv9hqgGxaWaWfLWe0
f5VmMdTGBTap9R3TnH6UOl1O8UeZ5Sdmlb1gF9eWtwRCoFFqq1qGH725eVtz7SazMqhc+iAAzCqg
l3cz4UajoST1fj6HD2Vfji5JOOL9COJ0HB1tfKk+Iv42GdE7CR3mOeWwiIctSa2oFETqcy8JeXIR
pQVjeJptd+ncdx22crPyt6lSOgQskXknCY0Wtqab2q52KMYdKLfwlQrCgmv0IvjfkSOgL2jmP6fZ
kWwt619DkGCfp6joqlt5cPIp2ya1hvm/zhjfLRB75DxksYbCMZ5JCHbtt+eUKEbZxUmRKlbxBY6D
ZByiFpU+3tpj0ChGLeCi2fu3ptz0N64H3Au5pCTj8fp88ZtR9c+UYe8OEh6u1x2TTyFGeyEvKVSA
zFqD/4MUe0iSfEBoJ5gN4uirx1XexEonkSdujQfNWMmSrYRvFu0Mtfd+5dlhnQvdKpZ40nYMgowf
0WuWa1T+Fh0MZVrGFOBMw0Gcljz478WA09bgbnh8m10RvWAeJXHbJyqrePdtZl0UhINIpsay/56F
MOHNqlDMmJIHs752AnJ3VHIc4J48pqXiO+Hb1L9+hTXG+NhXZ1/+eYdpyuUeMcrF4N4dhyr0gFNO
+ZRS6RvC9nFm9N0ZmMDROWqQAvT+pipzrjtUMHdsMlCzxSx/b6TbcQEfPrC/lj5K1XNBLlRRvGBP
C9qb3124hPiDaW0sUMqE8PwRnCNqx2kwUhyq2d97W1AXbTOUkMGvwxy7TsMGj1JrOo/FSFkxpVGE
uGUjhp3saaUOXZ8P4ehGrX2bZq7H6TSRn0IHx+8K1iEBQx4vItkLB0D/pnEvbMEPoepsTisIu8yg
GyJuzSacO5+C4y2xBwyUjRBU6T9RR3d1J5qkORGkn4BQPcgv0CB9vf3qXuIJ83YifbjkJ9W259OP
mbYjpnUL//tQ+mxJYCLu6riXaS4QUwQa4xxYY/y59Q1G+p4pnG5oXUZCLFDny2Y8FX0dRGsIHxbk
OgchJC18R9OSTUcdmP3iDuWFu2ccegQ+FSqyCIZYzrOGS8wx6G0SsIs/OQKab07LROa4foXL9jx4
55w83Ujt4Pmzjv42pJkrQejbEUtJYCCb/Uwqz+VheoW/H81LvwZUo+xnc/Gmk68FXGOipZtj7n05
+j4LblfV5wo7MY4R1m42OGPQniuofk3PsruwUIuN0j53A0i7YvuigTjoeon+9TBFxDnsVy+sTVH/
wNWW948A6jGJH2WyLiEgP9WHL9QDJ+aCXBQNsw1k5yitrWflRWfHWi9YHBif7nLokWyNAd3vAJkK
V90nFz9O7CMCPAlI/48aFbUXiTNotMk8GwJ9AVIsPmh+cxT6Ej8qJmXTIqQ2w9ty46SCyKCbpQjF
nPFD5K+uE/3b9J8X73X69WWnyJoKWTro+1SqpO28G65B4XFhTgYwh9WnuqY/xJXu5h7R5XKUyPq5
6nHfS1ZhZ15AARTwjDlc7xELOoYrB7NA8UrP1FLs5P2uItndjOcoBkT+SOpBIdGjev5DWW4f2t7t
SC4Yh/1FuMUBBdp2EZ4Y2ezu/+BHnrnOchJBCFGh1h59B78S9iLk86io+Pp+3M+B7Tn25DFZjbDd
D6WHNsHybaUfFDXuYNVnCctdnGrBAyuFTYo+t/wjzvVD/IFnavBpszBqr9tK7GfipSMM0HfawHOs
zwHyTKCDyss8xSXUEwSBmruaH8MVkz6veEpJBiGx2jBE0TFHZ6TBsVax0hhQ3zgosD38rAUwBNMf
VfRaVHCY/OFjXEdhd/+OoaZHD3gsLt7/Kp41fbfiGQ3vctt2/6ZTtlMQx6bc/3gn6sBGGa908Y0m
FWsxJFv8gr8hHH0Iy0rZfdhyfQBwfyafnXyYDUDtX3GXT7KIHf4ZxhdL27bUYrz7S3z8XVquFgEZ
sq6KsD27emuxzFHxRzBdoM1em8X2Q4c5uBDhHfLcTqn2YodxcHCFWQgOl4IEXDWvEWjgBq2KpUxg
hzIhc4gVvVgVCqYOpvqEfudhgWlk5fleLKaj6D5CJCisRzsOLM4qIc+pgcfNp4QJqAmaD18xEmzh
u8qcD/g9I9yfzx9hNVy9bnBFLO4YBN+PXn/UbgThyTnvgg2tFOrHCwAK0nkY7W1HLhTu9/923s/V
92LuBPAtNFoIRjXNoMq0JozEYmgq6ycIjDi7ZSJnQf9cE2Yd63/HhfSEQSiCaMZdkvAbardGoQMU
iN11tMDU3jxQQgfc0Odf4N6RTn0NqE1bKrUX8ciZGPllmgXnIxuXUKTMZXiA0lYVLfy86paKaNzu
Tjl2DJn6itcCV4t72QgJ+yj65Cwf4rRMkPphy7mHEgUS4CqSfm8v4QTUIxrRMFTOzCBFJ2tB65oz
nD7fAGD+/yIMG+sl7qwh2cevKeY3ZUlJWZGEKN1SZRtKRzKL8XOoY6HaTaTjWhC5B5Te1BEW2143
994VQ7Ji/h8a+bpj1s4c6X1LmLoQOj0xRq/uuu/1ciGOgCNTz+Bl/G7QWl7qgL0H0oNAkLhq8gr5
qTBkWGUh4/3Ay2W7+y1cPV85k44Ew/ksKCll50XtpqV+Ds49kHOfVh/C2fTJjWq7QOVWIRMr6VcF
rSLnXiQddxxndAg1RdutxAFDkr4R2PSicZKNReEX5D/YJOhqyI6eklfA9VW9+/mnHpLp0WkfYS7L
GEWGfYl117wt319bFoWRpB9lNySUJpXpcFswgbLgMjQJWFBBM6MKhMFCIgvA35bDYKTsG06tIZtx
jM9/9vuzR2edkXMR01aoYca9NemGY7IVOjpjMtvabG+vwqQNAMmcr0f6WD0jWB+nYGWIBsALSzBz
D2LEmHtkDDB2ECk7TuWsgl/UzkKgi5V+OUtE6ubah0pCMPQH+Y2US2ulotPmg6Uy+PgAP0KiygsC
gKxqvgSy4uisvFAkhgXI9VvXD1CMfFsjcXQJmKhgfR5cGfMg+I1J/TUHvtLpEnuzYeUVT1PfdW1L
+SKx2rpb3891EgD+baOvqUjLXZSoCqS3CUsoOCRG27sXL456HdOiD68oyT4ETyPnxl4XRg9zwpYi
S2bvKsQAgQDDqPwcwZAVEYKLSohP0gUgS/WMK2JM/+nWBHeIukDlWDNC3TPpE/JAFsqONMdMNVvS
fWAHre19a6hHCkKpPgg4Ir8l2a9JguycE/HxPJyQMPyUn4jqEfbhMzQ7BFM0lyhvnCThaFwCXabX
MmQ9Ss4+OMhxtkveu06EtKz64rfgiTRZXwSXr2aaka1j1C7DQGeL1mE8RQc2teTxY+TU7ge+y8oW
MVqaEHgIModeKW1zt+fQpSicrRDvCvE05G54ixuFurraUPFhrYJorsbW12JlF43h8OFXGyAj075/
4b7W28YXI6pZyLKFbIfT/iIpvgATBF6LEuFHvMPMr91xg+JvWckWtzLhk0YFPElYh2JoqY14Jgqy
FszKe82D7GUA6oEkGmA2of/7rXxVhCDOgjXKaZQMCYTfba8Xo/SntNr8tTqYFatPw4Qa+dyBOa3k
hzOT97jyqJ9X49vXtRK3BeLBfPOLt3fatAv4A1SRTM5ex+s3+irqKDqRuT9DUF/djQeZKWJNqzjU
Kby8M8Y/0terQEGBGQc3By/sl3DDeyYigBiajkiSe/Vi1qQqYlvGbAW2WAr76mIs4dSV7cd6+Azm
g2P38b1Nh5ivmPYIs0HhnU4uVvD7QLaynXMILIR/WaL2kcXvTC2OfN2WklW1UiHmFArHHy9hpr7M
F6FrloUMFJukhYrWx1WB6DO4b+RdFpPZrhyrNxMIBtFBSaxUNe8pRGkTEyMnV3dX9GLjIgIK4hVk
k9ZkeCFcZr01/09SKZhHElmQTsWKh6hbXWjEhiIRvPnXxpI5TylH8BoIq1hIYI37GA27ig4gVPLZ
kVQZFh/Vbn+eQXfneI3p1/rmFSi/JJ1a9WTWv+L2muOHzXC6zjR8x4Wm0rpWBNC72frwoTFL5AVl
hkzGtp4TMALh2gVnWCtx9tPhD9deA3R+AyGB1RJNPGn9jGl+gViCUljWw/XJ+uBnPLut8UZI4lIJ
SVK6m3zz/aYbeWuk3qFYlm77ULp7m6HAKNCUZ3d3IlvmEseHrWSHLESVHyW3HKAlVIMqJA3KgpZa
SZcW4WeDPvXO7a1sY/JM1nHmMpdXSbNqhOC7lFA2U2fwZ5y+N37Ah0Q1yAKCGt0LMVq3hW8k0ILm
6nbTY9Ag76H6f1fkjbGIQKUMYJSo6bB5mdHY4ZGLCpCgvZ9CUIlWjM7LQkcvrYyJdvI6rb9cX/G0
KkzS1Q8DnaL5X+5RG22D1UbXVHn5C3JKI4JiKEiXO7ELiSDo+6tZr5ckF592N/7gc7GFbXPJxvfF
gFxscw81pRgABuqA21uZ6W5mjdcAf+aFfdv4yLoCUgkqtuyIjQ7FrnzeQ495a8+J6GlBzNfLwlsP
KKvmbrxVtIkM7wJjKzp85hZtBKJhU1YwXJ5zS30fD9gAr0QcAd/rPQt1BW1P+N1kDdhy1cPlxTYN
uyqjuKPMQyNqNGnEXzYDTZQwOCUmUO1c7kn/3Xu8Po55a2UhnYzkzn6gn9QCvXquVjp9yr2YnvmZ
TkQXlaV9j2snAbuWDgIDopvKwzqRSlWdzx8IiJvNZ6DeMRAg4Wfphw3QGfGYdfF+iEPg/qraCQsR
jzOFlF1uYezHcAas6Xd9lbLICBrbxXdfPNXRDT0Xgqj7Z6S9FB9EQ9hnd5UXuGtqGpdKlgw7Z6PU
gMkWspWt3cBNtAL2Q0554DgY9qAge6YTpgO2XvpG3tBt6STBmlWfPt0+RrHhyiUP1NVHu24HJg+b
Dx4vF0C06ry8TB9t0+edqlTSWZ3QcVRU/gQOG6WRNS64uQ3z3x5+++heogvizErLy9aDd2l0/Zol
TJgXAsH+u1S4sem4E5sKjDofKuYCsgNhN+pJ7/R9gPRHUcDIrJ5WxjuGi09J/KeCYoKbHHurzobf
5sa33ZFD4vjiCGPJxi4fZAs62tgH4Lb9WRNs/E0eWsVlncA4hs9U8kLGLlbRmta3yYGMQPHUtBco
PLIrwZ8UoLmpX4WgpJZSsfbAeq25P5/iKZWHEEfkAzBjphw3BCj26Xl06B7Q0tTfe10j3AoH7LfU
9bM8gcXSOK2m2XlSDtlul0uzWmNHSbVLvclVP8FmNtDi512khebNJXuIVwEg7N6hCflybZ4INTyH
ifwMHNgbu9JjXGdU3Y2HkmnlZkU4nRu5hb9ntbsx3HrRIWpO7WqAlZtSmLhRZX4FxIp0/+oCJqmf
KY8fmJ8P3xOvHSIIxLQruE1HoK6scwdi1CMOoaI77wBRavdG5XxxLs7SKBtOwfWsFcO5kRJsCj+r
fadsXFRtxfsL0uKlZdyZuXUaKR0jNqoKc5Xg0Gle9KhsAORBRMz/Z7bG0jyNaqIzjPE/h9pfZ0K1
oRZkBsNQNWNqG+nm/mPU+DDYHJey0dPrwrROd1uuT04FZiLk9uSWptoBMJ/hpwm8eDfY6W49Bbqg
E/MEB0h/WiHQE36wsGEWnp1itXjBXscRpyehcKWv85cf1sasGxwZKUDHDoIlAoZ7yQFqyFItnJi5
gFDpp2pEJBlTs6h+ixD4wwgvvoDqoJd3+ZXHZq7kVl1tOG96nrpSDXn5Yvfqt9G+nKn2AGxnZMju
nIj+Qocr4OStqzDyAXArJHcQEUs3Ae/8FXhYIL4nUu687D5NhVrieu560I73tYfCu0c5mavjX8yZ
Lyzs2pHFBrsxBmBN5Nwp4klWpW7q4BJydKRKXO0NX900ZjDpzb87L1TYI/Zg1y/LOYuJF3o5APm8
F7I85Ir5OlOlCTEjVDBJI/EDmPMQZZwbOwF8FH5dLmp7bu6ln539qOj5Lo0YagqggGhLp001Pzgx
geQFQkoU8DolXTXBQGqfxNjxie6xy3ybzrkW3NPsr8zhh58/nb9gbKlZAt8EvGadUZFLI9RkI1uo
26Ty6SVX7tzLeHF4Mq78HDq1Vb/sLHXzEtCc9de0V5OCCpxbTZKZ5qPJql8MEae18OknXlHThoaP
fCIuPdaG06ECnd4LVz7S4hbjMSkI+1WzBWP+JHZOjlfwJMA43vwzi4M0v9dlouZeIdwQzX0onQo/
bVwSuhlgccPtcMtArSvDQn9C8gNVPQJVSUAPER4+HEIKFV+BqES7AMcuPKXgB0DtQJK7799cwpHq
zginJRXwzP8BhbYeeiWt4Iw8K71zNutFm9SSnFSTEsTcQ7gLi3OFtRHj8rr03AsokkPQI7fc/g14
MgbCa2jnEarm5fXanDzCBzfeuzJ/FonlfOorjFACjUYEUUXu3xsGzdjGt+8IapYZ2lU6LXeFRQpy
m7wAIv3KHxrDX7n+feL7OEk/UVtmh4pidNffgZFQ186j676wttLBIpH1zrAB+aIwIP896AUMdpZv
DoziBFqxe7xnDIiVGGuul4vzDIoaAhL/kDvAQZGEAtLjFtVZJFWtWPH1EH77LHTpl+jE9PThctul
ZUKi9IDyYHcNadbN8JvTEwMEtsETh7tEA5//YlzHxZ/uESTGAxp+bmLo4gMgaklsynf3b+VyNOrg
Yx2ihtskb6WOtSZJBgycdpcP08tIiI3alFReH21DzsTBC+rcc4gh3HnJUFoZ65g35G8tI0HS+p8C
BNMNMBju/s+mxtusViW2xEzBJ7cMnUiZw+G4a5KebJNSDyQhkWsN7NVoI15a0Vuw9A6p0Zgi9AtL
1nt74W8wGgprDJK71mPWEILlV8nW9WwTWMxqajmhCt12RZoyVgQ1KC9vV5wZgAQuZGTUiGWllwv2
yJruqQkK8rOm5/uPst3Tw9Xo37mS2A2dD7Rx7jX9g5h0a+vB7DuuoLD3g/glmK3v116OovzyJZyj
KMsRpGPw/emx1qhYLmk40zDOD8P/RkZQJxMZijGZsNkGMJYCfp6bdjJ+KoaiUcK3jgZdIGpI7BM5
hc6Q3vpu//05YHwYkV+XfAdFc+/P55aYVQJa2ExFehdZ5Hdv+X0XFDesm9YvqOwqGi5WR9wPUK9+
C6oR0gZruXLM+cUoolQZaZtpKHYUa11+cX0b0fflcyq1D/0jZyXSMQMGqp5crh7e/9I5IPVP7qrU
sUbjCiFGixaSEhzQpJWjSIixBKQpEwYQFAxIFgNueVVzuFSYUd1hZJKQqjccTgsXx47mPh/YFFEL
T/UbVOytOD8eMhEBRj9Pq+nfwSCzPgxqOk1YdOOnuhfbUDDw3UEoddG8XooOVDew7h1VAgznCmZb
bWL0I6AuVwEzNo+2eA4SV0RuWngIYxmzlaRX1jdA6GHUIEkuekvJhSqiCt5ENb1uHf+iBGWip87x
yTpeWlX8+InqRyQkTKpJtie5x0ajQVh+lG5IgjuGTYS0hFlQ2qUvETqAfOOcppYks8cjbLO48rUD
227P2HWmliu8bVh3b1hqzSB+2IdVXi/97UZ4SbHRJKyEAXU/fzcWB2zKWsmuS0di5Z3t6TbWwDNZ
bCV5szD3g4zwbxW0oF+EZnNite/+pN8AaMG8lzzT7M6t6+8KHHAF2VT+xLiWHG//qqbN7tBignOv
r7oobHqAMLXDNqdm4gqg7RMO3JORGQzCJLy4exnHcBTLUDhSFKas9F3DnDDk9/+/V7ks9V4iWP5i
H6bcM7lvTtbRpx+Cfe92/3eoYuZUjRvli7JubxJ6C8IJ+1LpIijlEyxND09ubDzlbExjnES1tzFz
hU4WAbLifC8sPMOE8l7cB2QKalJHpuIjHNAZkmX/Mtu8nykPy2sTrn+tf9aFmfZSedumCTCKI8/1
75JFRqu447YMWUIkguFtXD5i/VcTo9jBenhslX1bh6WmESZOJgPbkZ1sRIgr4vKtgJBFu0Cr1c22
2ClTdZJdl9MME62sis241+IeO5pRxCnPXF9yh/4OoQHRKoHSaTLGiEl0OgIrHwZHdFE8VK57ZuS2
cyjLKuci/rhEV2liu6Ez46nS6wBxg9zU/WehfS/rJbSIfE1bNa3zcMCv9u9B9OFfKI9yPWooqO1Y
W+/ySTzuumMxu/VbIa2SY8BnriEv+C6GsX4DImaV0W38nX1CK/Y8EmUEvpcF89W6wKBmAHKVRKZ5
nrMrXyhTg3ZBpwlJQSzjhBnlSpShWJqsQjpF0S258OjJe8cqbCAPvYnVgI+S3zqW0YjgSVFPGdue
Ix5akrcJ0Tm318dvGyQKcF21NExodDGJOw8GHHo2ajRCxf/1N3yL9/MGq9UX8ms1MNccs76dvTbH
FOQWEjK/IdquA9yRArRoVrqYene7iLM2g8rKbhvUDc+XHv0Sx/mPv7Pj/cYzUNJITwuBedv+FaqL
j5cwDk67K6UW3XLvqrZGp1YdpUrNiArJxLdbPCkcc2grBesNk+z1wvOPK/jhs3MY49x4nwsFQHAt
sS9lCbUqAZgIATM4kT1nztnlxQ3pjWiNgum3KwxR3Z8UHbqaRSAh33jiqbF9BCGM6Fv4drd4BD9L
s6LjODY2utx8sEz+lMGtU1gB4b7brVI2KW6TBhyJK76F0s7vSKsGlyg5/bQe/83o+N1uS0yBtWe9
plOFzm16RTkhRto/eWKxp4pvVa5GLWvAzNd+OQpsy4YQe+w3b/7TmKv4+elcD9+SOHt2C+dqUS5n
jsrbH2LLq6qt6x+mZgV/+iTr1FEOpNVJwnc0IVoXIc0pHe5Rjj2A0pawAYvqf8z32RQOUQZ5CVPa
EbRlA8RCAVlF0cinT/9wd2M4TDOdEY2mWdmIC7jQ6AOHg/6ti77imDrzUBbcTnFAKU/4mysKnSpQ
Z0F2nEeaROUu3SrMCAJcDEfDwNKtnaz+YCacCV1354Jt2iH7qh0xacNfI0aB/O+KmTiuC79m8KlA
tQnfNYu/OttpdkXJ6XQxl5lPxa7HX+eklZwp0Lb82QdIgGwkcGIwAWK65ZpRyTzdLu0yegt99BeD
XH483ZvdeDCJExKLak8Hs30oHYtYb3pL1jSNP96B2ahzO+4n3xtS8AUy733pi3Cf6JfDvmIIYG5Z
edFBZ/RMbck10Fmro9PHV94NflAR6EyoSdn/Z2dUk94Qnbn8w2zHiuvlgbYHPBFRxlbOZsndRNEq
hLDvL9+iO3CDmpJ11QhzsKwzZi2TVy5PXpV/HWf0uDSVr2iYvB+qy1KiVNVVpSBjb+7Ui1H030is
PgYUULjNYNC0aDxcEJ4Xgso2+iRM27LDMHmgiDtgVLq+R6+LndGsE1QwIBh3C+CCE3eB2hZ3v2wp
3UuS4pJ1Ixyyy+VJPz7kIzDlYZvoY4Ztki8suWojuV7vBaFd93LF7bALnFBTRPWs2wDOdj3YqDx+
DQ3AXbfwsP24SOjFjaNksZmkYd1JeT/RbqxuoxWfz0TnOmtLPdUZR+4shGbAzexZc1iGrJB63gXT
sha1+Zxp2crt6mjAJoLEGjfBJ3Wyq3f1CkOHVFdXi+IHhnr6PGlGPuZjaEwWDDISpNSwRiWA0ooC
hIJnN3cJ78XXrBxfo3/IUl4ABFlrCOQWOCKJ2PTI2ASz6k1uUQh35XxxcYWdW9zmxji+1pTR/vfn
oNU/r9L4tdmgm8HwKMWfLVsPeul5WXCgLa5QdFyReyVfbVQ8KJd9HX1mAu6y6qowSljxDe7LX9/1
xWFhZ4ai10rUeS7FFXHQ9QD9OHijHfB+bhjaCZNCejnz/7wX1ITrA/ZTx4Ds4H+dunZoIlc9cioL
hfVkGWEIOeNhmrxtqXzTeORbCWLdnsUWbSwuh3yxKJwtrpWqU0858ruuS7z00NIENJXxpFkyVSlb
i2l05wWarz2VBswX8GeKcp6HZXPegituUj6oG4nUq81gJF9qAoFhav5/WgXcGjXpV6R+eqd7sQP7
ayzowMRs+5RpXaFjhq+TSijBfRK6WfC5jus7zy9gknliMNH8P8kZH1BPDRwdyz9K68X59/FQBcyd
l0DcK56NX8DPqc3+QH/bMCHdU9DV8BcKGuD+AvmaS/OgdjVR9stpt3iQWW/iqgUnJZIsyDevjm+k
HsEcGiAra1mgLNB7Uk+J6SfufTlscTb5N7WLfABGKt/g74bTINiq9K82I/7YSkAH/8IDntau7UCT
BPxUyDOzW/yDF04Hntmse97hAdz6NPY0OesOY6ZdnVpzyyttJvYQS8d/H//w4A3EdhsCns8wLUiR
l51LzynAjzDP3cq/IgncmvC7O0uUWppKef97Aec4TIKGR45Mb0D3C2tY3z0bSRph0CSuePxod5TR
lffEJvbxuCVO0gVjyx5tipI/4mFFfBmF/IjMHrzaMoCE0GpCAvjkJIIqReqg6yY4Wdwg/uu8Ke+U
2GP6w/75I96B2QHO9AkrJ9vp3GShZpd8y/bvlVE/HZlLr4VzDaZTAwuUIJqBgCBaiSQxIcheUywl
Q2wG1HXRNu91ksiEJbg4sz17gTBxNf4+wpyRkZ4ldl0N5jO+L/eHloCTjPN9NY3VkodSpMNuCgfT
6K9W1NjK53l4jL0qwf7TWp5HA1DKrpUz8/WNnct3eUF2Tjz7fcf212AQnB/stX2CfpNwPu9JbXYa
mE+JajjibLc00EnmxAni9JFzpgTnYbO7jAOh58ofj4ANQG1CrI7Jv1ZIV8hU1wFI9zRU9JL23FLK
0sixzQfNlrl58MGGxMi+gpO/5ik5Y4AmTXSAI0kfYo+atpRoSGNXCyxjxxtHX3ZnQuOo/k351w6V
BO77d562sNOw+COzkz04qDB+7ma+qpn8MR4M6Q0bh6ONUDQTHJ691jeAW8gTlYO8xmCvA2CtOwcT
fQ5+pbEsewD/ZfsRrZG4p59L2WbcbMcLRXWpnRc+3AI0mMI7eLsRv9WUjUteVrBNNUV+bAiknipr
dxoCDVDpUTXV1GDCZGb7q8vJ29AGR8OMxeA6M7R9bFmboaXrttCtodFzn3o/01HHJ1XHeDrYwloX
shog8kc1xPAT2yzlE9j8+vf0ut3RCVBKnIFv6JFHVjcNMfAuj7fFSBvBtiTcmeYkcVTV2iK4FZxP
WSU4vwD4KM2jp+zja5uqEzi+Z/XAUo1LNnCAD63316rGBBFM5WRIbOfVtXNjK6eSxF7l1ZOYOKIw
vfNNjXYLX6CbIL+ao5Pr/Q8kYjCSO1LLaK+x0TXFVqphtoXj+gKxAwJ7bMdEllICkJqJO7X+i0EE
zQu//CWmXYnXdgT1NM4gMEwzd2Ab87iTBgKqip6KePJN1u9fHsuNXjA4zc6y5Ej8g8fguz4SvS9/
HWZ98Pt9BOpnhEtLfDfdR2EetBhmvna2lnjt6Wg8v8RqbY9wFmDnC50eV2E3Wsr4IO8sYwhjyueH
W13asISfxRIb3StvZJNWReaboCuEnEbLPnXdb+FJC1k1SVAMhHa3paqp1PFr3xnrHh06mtZj6cr8
q6DMHdpbQ/Yx3b+1VNwuHkTOmih5S1FCXYAUkjDZir9T3ZrxxSjFXAt57+sN6c1fJ2XpLyMHR4tb
XsvrK1am1MplAJ0CQTU4Gc8dG/Jdddw0QKI7A8L8O4xg85PYDjT3UwYozlajbw+ldrnCSgHHFGal
wh1PJT9t/OOniQNLKtiS20ArDlRa4lMtyyvNrDgyBK0qrooV32zYwl+60ESA0aj/I6Gj5rELDIfl
GsZuZLocVCGej2XJrGpIL6ep3nkYmf47CWr2wHUFiBCdZE6KW2IwNJxc1WBkFx4JYXjw4MxhN+rn
wSJ+DNvh7HwSfRK1X8HnM6RIi+5fJ0p8x8X5LJUJ6Rj3VkZJhyNmK0A9Tp8Y+Lz9ArDislkDFcgU
h/TH0YeL0mqHGIptt6dUuY1aCIhFdRW4OPVEwtMrKtSv0zxYVwksNEuXGH8jDc/8n5lZRJFIEctr
gjQ0TjkmXPJJcaKMSKHl2fUNqQHNxZLpN4NGk0MOUGlMeRa4Q1OvTxPFatRm9iOTldKsr2QSP6oE
5dKAvxKO+1IpT9vqHVvZ+sAx7XGBd8cjmucDneOjs4b+RdycolFVvXJQAFXlOjma/EP79nni/EcD
lClTOUWQCyS+zq+X2+g31hxtfnxs+OtuGpnm/Re9qrNZ4jL2DQp0l2RkT22P6A0bzXGFRnhay7js
fguPoG8S+AunUFScJ1umW+CiCAiWO04qBGlmElVoZmeyFSJPv8lTGFZiyOkwFdXoGlIhY8EQJT8f
ACdpGyvcr9Kzps0+nnvlNtYjg9A+l2QkjkWmZRSFtI1nJVDWss7Tjmbl/VeOU30carTuEWQr6c3N
53BQ5n2dS9LZAFD/buc6SI6V8M/vCZFTAOiwWR5CJJuElMG57daF59WeIdRYBJ5M4QptxTEAJj5Y
koH4b1+AOlIsXygBKk+7jDaiBREEqjfC21OR9VTM/B0ZAbqciNvSxWh/ZL1yddqBD7jhd+Yh61Il
dSfgV1C+zrvm4xUbeRnaPUzOY0lZAGGqBl2dbroOTwzhybjDpfr7V68LWSFBnE2P+9pQ4diXIaZd
URZi8FVi2v5Pgi3xOaKre+eHfulpwdDQdWBK4WKnOwYcxybU85IpOM+RrklviTlpxwMRiqvdVJNw
THF9rhVbN3BsnlPbtNciF3oeQDHSPaiKTgbZsmkyZZWm9KfLmqk5XfLm8fHFUmnrzK7RWK572Yt5
oo1NqDH0sHDFw+oUXrX7IknRkZmWo1cjjA82CN0BU0GUrJM+KDvPvNcAMIHCbZXLoDAWnbUS+CFj
XLMJYazH7NlfhvlOHzEzuN9T3xNLAQNUoTLm0RUed0z5GA5KUkP/UDex+HOkaXhrdvTLT0TcH/mR
q7jCP6x1UrBr28MT11GXUOjLX0WkN8Jy065YaJOkMiUUFAGG7rFI2bL42mx3vTq/JaqLo5JPEdvE
AEVztOCx8bNJ1Jdn2CsM3VbYS9xqEhGQCkgm2cOa5B2HxdGhYl/MQ80o/EzUumW7ZnzSdCxDghAt
EU2Iw1XI6oOI6bv0jo/ODNjdsZfsRWItiTjhYj79WyzY1d5nuMpXVvijweUJFxYoEkC/W2+itosu
QHZiLkXlH9nt7lQBQPPEyGin4+/iPARbdktv+LCcVijovlXQtcpMkCIS929JnzcHH/AA0kUuYIrO
h1CA/JuHF9bsWZQ2rlAm+E3bNuAZcqd5vAUe/BOyHyYKeQwVKqwKOKLmkPrUiQQpQQIgh0ffC90k
BMd5hfuc/o8/5n3vVoWRyAMs04oDTUtQZ3mJVejzGAffrKAlB7QG70cNqOyn3bCwUllhFBirO+Bj
d5KgE7Q8F2bIP2tktu0XgVvWmeSnOP9saMBOMQv4r4NVDVu1eg2sTKD3k69HHDefoFnkQTuwJZwP
0AMPG3NgBMfBdiAI5B5ZSywCySaeQrF1vkIvJgngS21Os3s2Iom5GZTBXtJ3WmZszwWhbBUufzIZ
yqjUV2BLZ6oAboW82t0qpGTYYDAWUV0N/IHjo+pb7RCY3nFLd3n80darzkwoavIRUcEECndGN439
WZSM8IFzo8ASOPF1Cra8znWOh71/dK0vviby+MdJaOya9P1vUutZLQ2FBjWywNnGoiPGWXkslXmq
2j12b6t59kTaAwjRlF+q1yDUc6KyOiWgW9XMUpNT2giwJfL6hFDq3LpQrEcz8ptP5bC/8t1zXT//
UYM7xWcnUnC6Tu/za8sPL09eOfCaX8soZahqlkrRdWyQ62LSxXz3xLUQ1MyWI3MSES3nnjxlnIP2
Z4xEVVj065ekx7RhtsredTSmn7u0WiDEXMvf9J9xR9JvmwKjqSmksunHunsydbunh/doqYPh8hG8
J//4JHRZoiZCQW01/vSFdUrDkllebR0NGUWURuq/JTEBncvHRjTgSOHwi/0pOjiVMf3mM07DYgts
jVnST34NfhZYLTi3Dny7G9fog+ceMY0b6lBfg1DvCdDcjd18c/aJBO/M26XZiT6E1nTQxSt2iacp
p/Eb8GGBjj9R3W0yZ1CZeSSfmlqXb/vWVfGi40HGk21n5W6D8J8TnUv5ijzJtMs2r1UCM0t8YF++
DbnWn+WhPyJ5jTQuNq3uQlZfZ2+MjeJhRzcgB3FjtrdKZDxZxX7YSuP1iG3FC+NWuebGtsoVoQ0x
QCVKHN+jntQ/HEvWqIR8IgrULTkp7BPAcPG/ZSJAWIwSxjKcuQnz3eUD29FK80bUadempYfO8AkG
EQyTbUaNLWz2ayM9dF+30xlDCll4NVSrzz8ylnBD23a0v5tVbQRVOeM46usTz0SiLcN/VUqznP/I
F+V6D4RsuUiY9RVFMbUpJ7vdsXp2Q8HwQ7XWZpnun/oLDa9tH+7ZascboUw23DWv6ZO57xjbf0Sr
0HyNgHMi5Gpszgujga5dLZEYLA50jKYdqQw7IqPThXpB34JuPSJ+QFapI5wojVvIlYX/+YKCWzIb
ZmGT066ZGZWkxW7mjhpmHEifT/wbssBZxYzctJGqLbGMLCxL+LxT1lIetd9sp2cW2G1pH64oWoCU
Hz9VqbCgKssh6kMmDdxqluZx8MHjRoSR2ilkxxBR/QEcm1bBBJAhELWcboDGo5GuSn5lIyrliM9v
sKzKiGs/Zt94yIGO6WhfPJNCV5RTDXHYuvSPVOwUZwKPELFP6ANUamSqidEpYE0uZqCo0orDFrAd
vDy8lJJLY6BMu9zGiITcQTNQDicaUqjnw1JedhelgMtt5ytgxgfklY05lLnoN6QrJjaFLEzLMo71
5CWL+mkklev9x2LjA1zq/RLabv2BKldienK0TXHden0DL/r3XY0dwWbgUxLAQkbS3EJqSObEOpXo
j+gEJLYPCpelpxcj0MLOHSG4quSrB/qNspGzCO3CSp3Mm+VqB5ImNvc2kgLRc56Nt65rjPV9/jUX
cPzBmS5Pm9lllgtmP+GoADahYgRe8QxA+Wbj/mvP3oD5OUFpADofcwifgOA93xJMrjOOIuDqNAY7
Lz8hfzJHMb8AFr9UIAND6As8XNcHCJ3YoQhcREeQtRNRAxSV8O/KoVnBIi2fOheW4FO1qD+WQMif
P+/DSeyPxWtWY9wJCcUr5kYFG+KIgz2BMe9gMTwVjEQt/5iPInRQReBkzbQpE+AFNQaKseKABXci
AYRIwzLL+cV+kb85OV319uEOg+1iZ2XDQKv3rEvx1WZTguL7n0oDaqphkPJBthF4lOZgXKW11iX8
7+xeoqi3U2j0uv3K2cJlsgTc78yQP5FfaIzMBXhbbxvWzYMvPGGU6atpvW+f3g1fcw4LixWu1AuB
uNcNw5HrHboXsi4ra6B5I0OwQJXvKjcNN0aTTXqc9pEL/0G24GyE2F0kCaboWBIR8Q/+0Oz5gNg1
eXDj6E8S8ti8nPWiPal6p5tOGln8TZp454nTms/HaXcQW9VHDomTlQQboYLfZLu0GHYlBdhWBZoD
Jhl4m/NGTdRvCXzWSLZE/mjDDNf2g7IQPUMa7t4fFIMHNgBUbncUigvOpWWDvQmspB1qqyU9ANUf
M65PvTK9kqVQCL8nNrI9qHeAL3hpz6ckC/kxoPFqNtB4eZJow1Ozt7itCwdylwGE9MaV6MyP/qUc
XRKhRuoj93bwFjs89KV8E9ZdhIO8LYrGlvWPTcQbvKZBHtn84J9txozAFSx0BV+Djc5UNP1fWltl
36UsMwa7J0hgPqPjK3ATUARj3NO1wtsMCQidKFBrCCBwA8FS1ptzwPAhcnW+CmchD0dkGmslPwHs
PFqz1Ya1ILN+0nZvoJihdLKC4f5frflff3qILutkvizmzqLcWJNnoxoD1MHzdgUNbBoV0C7syVIQ
Q6bwPhAixNqlOS79rktq3iv6X1fQnopuxo4VcIclu1ygvrpRI85OcJWJwec5ZgqjpZ1Wr5ntutLX
AS7rgGrxo3schhxJme63QEbPE4Y3q4mW7ByDU5XGfM2w7m3vwTmhVbqEaCgykWx5wd/9nkfgTHw2
/1nwBsCi++4L9r6FFX3Q46Uwuey3pmsmMU9g4gt35A1YuVIIE5BomV8OMds/DyYlF7DLIfW3YlLN
Q9VlsvGKlZnqRCGJfppH5uUb7mqh6N0EIpNrvlPEZAbaNqc9oEqtevH3BlJQcVO4UKklqneXK8es
o74ql0te0tSh8ntYkspbbBRcQrbFU/Ls78oCmT6HZ+p1qYWWnZAOc5Z2RA51cp3rnz4gzbxKBB2T
2EPgAPBlQv1PCvlS5QuAZz2H+LtvzdiH8VtVfVvnrqQW2tcg0X1HkdHpXcl6NDjXoygj/kdwQejh
RCGrzmDjZch/GE2Cs2NUFnoY4ZS9N8p1Wr3qlP4SysANgzKx2VA75eON5dK4nwINfWJHhPt0HgXb
GIpHoGNUsnzY6Pe3NuoDGLzB/KL7zeIoRj77fdWOYOq99mLz9YWeK5Qhg218MX/VLghJslouiqs3
NQZTdMN60HFi2SsL7UT6/o/oNPo/e7F4NKGb3G/X2UWgglRDZuCnqdBCuUWl0jQ1hz6lJMo2hgyW
D6gH4QSHcPjEaWDzrBmQZBXJwLJ614atpmqGGTf3rNjIku9Hib1Cn+yaMizYVXht4f6OmmYeRj1a
GovQVNOc5a8axoPUbbKtABPRfs+rQVjZF+UHKEKSAsHqIU8aS6/0xdP6UOV6ElZzUQpDxsiS3Nvi
LGRAGLFaGINSwkQQ9a0lI2DgNYm9SQS+ymIGfXvUUQKCuS8w2QbO1LL9t1OC7qcNXYSGlbHdOaJh
u46a5Ph+nfivM0jnwGiogwnmLwyPx0Bkg8gmmQ/mtAcaW69EtZ0yKIcAPh1Ky2SlIo92fWZ3anT/
P+y9tbR22CNAyHGOPZlz5/W35nVJ9MiiOHbKvoUt9SwlJwEC+/hqc7kCShn2vYZK0zijSCTw2GJa
c+x6SrGdjctkj3FXxL52E0K+xDjE2WIIRwYjgi0X+kS/s5Z2OqswdbP2k+EqvUYp0d++5E25yf28
zaI61Clk5PxpIDadk8WWDuVVyQoX6CINCO2gk+Y2XL1VVftq2sky5yn4IjzT4YkH9D7OXU93s6dR
Q6lxqoYvFENTvsjMWgDbMr8AX97xk143Tb+CL8htGgXUDUAOfyHjyU2mNHhov3dQYbjQIzKLea3o
pKg+Uxcuy96KQGOb+7Bs+TCipiVLpz0ilGBIQ8sBXZBaW7TlTFneEGDNe8vu6ZbkFsRelm8frUAs
1Ph8obZHPUcBlONpxkTbkCnADV4brJOpLd7w19qDtHCqDC9Xy1mBM6NZFOYm45j1Yd5d8sg/anPI
ArDPu3frqi8mLMdmF+zR2Zehx77vRIumVl9j2FcqdXyWJ6BrAjfnRQA4q64JUBbym3MjceF566wP
fqMdKSHO7Yrk/P1SyBr2IrWosn1z+04PV2L1+bCz2tsZ1md2aSnWft8FeR+ni7vpZHrmQUsfW4Bq
aMiwg028DXcVz/62NwSTekwGXNOVWjezTGZYFl1JjuFgJRZneE3bGXa4t3kRqdh2yW6FQu8/QEjf
xBZxoUhEVzVh1RBiwBE97hcx45SzTp7FBk7yJLEYG+GEIRc4Ef//G4Rs6Ilwz3FeOxYHjR0Arx2v
u+OBOv/Jjv+48ZPqXPWp2znqL132uQfDKfew948Bij9i/Slw/ywUnsPlm04WAHJmJ/rEZTZJOVvC
GSkiruAPVLcgaM1ldBPU5RW+KVqmCDBo+Ikmg5CeyCGLfo+9i1y23D8C9V7C3xW6NoLDwFe0GU26
aDcvVPLxEa7N555AtPqlu3vEkuDMXwaXC5B37HN3HD8wMlVD+QgcrlMqrgN3EnhRta4qNQP5Hy+R
XTBCxEGl7Yk8jifNwwzXj0dt92AqHWwC/9XvwVcIR3XH4LcG47xaBM5boP751/pD9jTzEN1I0LUW
KgyfF/NriYI9MzWGkRPrmlQyql5onuFiqrouo66XKuyT2tP0qV/84hh5c8LwalSSalJhOFakC6XH
Lj1wDl6UwGwdUiTWt9sU6EjEMDoJ26/rWoi0a28b1xFyk62gMPQDJXke7UYXxxg/rR2kGdHXiJwJ
pRG5CilmOxW3MWxsQlka6s9eAS3/j7OQbeh+xBK3KIKsDwtGikNOJEK0yVfLQy2HTL1k/Phe8/yi
grvBODSWOLfMRglD0GwB6xVfWcXzO0suyNct9dZL9iRP9nQLBAX1fF0JEvPzzsHbYprpCPRrL6tt
kf8Xb81aIqBnaS79E2HJvIc2YjJT95jXxkqD8K6zTuY4LsRVF8PSuHewvd3Fb75PHQ9uPNQuVt+U
lyug7sUJUeSeLgVhKoKkH7MlbhHXIPNtHS9svKqPeDOEAv2fRgfikDS0T9N+luZOwQLatjdqsrkb
JD4+QElFxIn55XKGniFH8WBEutEEGK/+qgejmOYBKc7jTGmSZN+UPCeiKT95gDnfIEhAWOs6tf4v
0wfBXnHS6ybEOteZg99uaKY4nCUE6kEATmdUWoESL/Z1GNzPsisp9b87eU+V0bZcjUu+BQ37oJf/
JW2MRJ2AQl2faoedWyLBrqA5dAW4EUrM6DUK0j4pMsJby0T2axuP3XseIToYTkt6DCkPQZX0ewOd
TJHQEhQXv0K4JF4sIMyzc0Sg2s3ElPRat6cFNOxb+G1wUuVRWCuvCWmpBV3ftF0FOgzPIe0Ko/Ia
LSKKlyWcKkdUzUV6DmJzIIXC8rF0v0SXaQCJE6FzQcCggWrVRMICesZYAu633Ca1k4XYzEoxAs+U
+X2sSsepzAM4pdqSyoznrWztZaiX9FbH42NTzq0fL3w94BkmVGfx0iDnfbAduS4KOyeVwo1Q44p6
PZXXCIYk/+zcr39CcYTY7j4c38NsPBC6mipdSRGBT8xliAamwaV5YrXjjvjXAKrv/TTGpLcPrqPD
1lF+Ll3HegClRTrV9C5NTVdUeY2RDK868iVgnAHWkcWdK/39/9nzNwUUuIjJZepsCetdfWwG/yBj
Ojiy+i/ADlwhN2tBR2k3IWNrDVYyR+rQFJ+KxR45nPy+8Pf+klNeaSOrQbOUBdQfvH1UToDTlVqw
UdnmZuB+bsay7yJFiLlOVE8HgN7qDOmvacHjamTI+oaEPxJTv8lyS4DmvAIo2CgdUE/UrvuHX8lc
OsKvAIoV2fP2v2VNSWF0ZElUSYYcIA7T1mtiWdmx8AX2+/ZBBOmwQYXiInWwQJtbSloCtTVCiciF
5WtQ7xQ1T2lLe7I+sScL0AktCnslvUcRXBevOCjD7FOJXvfKEZj83MNMtPKC89nGG5c0f+wSMlPd
YJFku7RBOovQQtqTgO8frZHzZkZuLFvNGe1Qo7lBQWmobwVr1THDvsEUzQ5dlOnv95+Gq/6e6moP
pGpFV+ce2EC71KuEOj98zqKat8OSeY5vvYvNghfAAC3kbKaOKer357uM4ZwUF7KcUvSl0JKXCIVf
ggyXVGkAQlE8uoO5YUag0OgZRTSN5Kz0MoYtXI6L4ssP9vhsZjKYao69L9jeN0V+W/wBA14axUM7
moYonFWS2ajuY7AOheXzSoG9uMXM2ERvcfd8Zn8QEFdnm0HEjKtT54RnoBSDKdlA/EA8cnG12xiX
jH7ATA/XsWqG2ZIgKxYm5PO4zQNhgjNpNE8cfYovv3yn6lWRSggmNlGce0/6pSmBvealVhHEBJTa
Lkw1MgeD3hSKhd2pu0A9a2x8AH+ktOyWW+TkB36Od+bLg8aHRyVa5CTijudPjmgud7Eaix97Tcks
yD9tLNw65YgQsjAGE9UKsDecAEjwyo8rNe9nNEIoyRIJ93SIYcVpIoYCp66glYq+WtbaU9N7is8A
1cY6o8FlgzJ/U5gm275w57MtqncXQZSljZn0UnqsHbpGXQCuNMit8uxm1sLD83BVoGMS7ROomOLS
+FOVERuXvn0lKRLcYGpr74ziNpABFbfZj40PMls9PWIf8p92NSGQxBsuijYNP3eJW2ZsFIit3qDW
HTtsi2m6azkJTpRA6qYrtFGpIRYbeoSkLPqSryMj/pdK0PwUD7w5AWJmx3dMaVF8KdhHpg7k36he
sKqNl56mpq5nEzN/WngnJql5blIPUu+KnDRXY5CTYf/2nrn9k2eqoa05AbG7+7iu/c8JhRC2d4e4
OGHP8P5geaWQGmwW5eyCMog5CcWZoxEHE8hhyvd2/yX354JCX2nowLkYszCpZlN4KLvbbm5a1t4j
j9CasPUwRNYWHPE7hPM/39UJX2bYyo9dasbnNnLworCaUF7M/8w3evtouXV2bmSaribzrfBSUxwf
2mecHB9V5c2sMRdPC1EdLVCfgL0cE7ET9A8CPYqVvB5Q8/kT3AOzEQYBFJNk26a1posgLY8G4+ts
Tft3X0o6+5dgGcld8BRgglYzXVg+1prbVYWAlf7tfC/JaTojJvAcnuSBRB0H9mjooWEoOcLivS43
17vRnndY04jb2gbLYq6pFs//IBOaAkpySQhGNHWsCYA+ojhnxJV4ceY5T++3I7ENDzjPCVbNEgWh
27e8Mh6PczOogmseOMXZdIpStUTnQJo22DVd5gImIQgmfZofjF4/NF1I9Rnpb++/PMnKIA67+DHK
P/0vhZKBoDFT1c7y/abHMo9rPznbsXvWAJjOk86Uyr8rd5zUaL/3dnXnthQXkwh36bGaVN1EpsXG
DjzpSkCU4oLDtKAjDSpB8IDUk7QHd2npZt16ulkTwouKppJJMVe8WQnAck299LO/jJyLK/mUdO6S
yFWtlqFGz3ciDiiTtpUXDTEOduFFM9f/+qHp0Z9xtYZ9Nlb6MuQ+s7KkvqiX24ID5Rlbt5q7frQo
xPSh8uJ458+TIx1ZzxR2XzvpziHCcSPDW4F1wxlyJfUbUpgdHt+n72gGUZOK7xGTrc9rQ5oJ7mmi
HgmMSMtzhvrSgcvZg2LSFaGk8uSC0hF/GaPZUMFFK7K/TUORDScZaDWmQBzUko3o8FP3C/gsU4jU
TPtWr53gONhBqqjqWMsRU2GrFbQruKs5wwZdsUOZ5hP6mL3BAPPQcJCYCNgQVIphgeeC/cEV9+1t
tBigxFOhSddsHqzLDzlDYhAc2QGbBVCENnmPDq9R2LM6I9bnfYxMK6KuaXrf72XUskrtz6c6aFGX
jsO9HRUEO0WuMs+XhDYNr8AUL5Bz9gzRxZWfeQMvx2zDwP1h0Qg4qj/cKK+UEbavTywQYt7TB8CC
r/Ek5KOSHUoNbPdU5x/gMEbtD7OB93dejVP7seWnI5PlOqPLC7u5jM5TFj7msL43nmqZ+Nzm5WCd
OY8e8VSGgzkyN11qqEOMzK54oZ+JNlWa8honED7JsrMpnQVXjyEJOW4uPty70bTOALJ94aSRtfeI
2uRobQNJMA+celzRGNsYEmHhCBF7iuYUmC7RYlGCCUZ97BWuCITnt3f0bnt+aRNlsHTJBN97/5qD
4AW5gZ4+h0nKEae2rDPoIXOWy3xGcvAk8mlSAT2nZ0e7slO+cOOtLYxAPMnfyr0yqytNhyImm/Tg
vfQj9zjckQIgYJ+lV0sj5xFWKycR1hUof7yii2IGWuaP7N6WAwl27K8DgccmoI3VA8EZTeWLjQh8
e7rMQWArWF0FnZSWVeRZdW87Dx7xYqNS9n0RcMvK0Hon7PNNJrp+/CYVq/z6G4M2Lk5zq4RR6NO6
y1gQilG5aSKG8IZ6K/G1ToyHRCs0nLA+e6RPtw3sstMsRT+E4PbSTRToYQvdH4nP8S0+93UdZB1J
gGPPsFlx/2H7XYJTtH0iUBHHgr5iQ0KoJWsiNbM8SYjwkIxbnQCJrwgctYCElQSsSu2PnkqM/ScL
ubSHYHbwRJ6wtNcdM02k/e7IrtGy+aUAD0Jr38nIrDxPxJzU64gAwpvJSuftsVumNKxuUdKpJ/Bd
75ZHrfDGIEW81GAYvmJk2wpth73FZnclyNpgtIrIv4yWvtwRwY/Ieu4ynAg1bPcBppKWUh3lxfNl
cx5Qn+kliIqzHq9pF+oJ+L+vYRG/RNLcPt5eSgH5ENbl+14GQMKjI6AhxJqdSkoQ1gEJc2bCvtmL
KYR8O5pvnt7Szj82JjNvAlDHM9GtI21xN2zNcjAzsm0ANAK8GzchqwpjQEEUu3Pn/8Qf+eZoHEWm
3QPQP76yG8+XT9diSYUM3rn9aR1gfV8swqSFx/a5KqO9g7spnuY/aoHKSkDtQpegholQ7qNHsO5J
vo3qWP4XwTrFVMM7uDyVtiPM75ElFFWFxmVlTCVwYq97ssJqrIDvR7gvRUvRaeckkCW5aUZDA8R+
rHxkz9uF4dPimOyXMG+yq9BffMzit5oIJzaqP+ddaixT4T+KXre4A22KC3qzQi9gtgZhy0+gkMuD
3weZmoWVv9kU/SWzP0mwAO89d0clU0mpLT5vmY4rJw+z7jDN5dQMMvpA7ts/N4tQ89dTgyXjM5Eq
jssYaZX55818TX0O5YeTvJm3mvoGoo6JLhvXBDg89GT25XXACJ2xVqgpi1c3CgHILGB2r23J5nxN
u3zAw8CD8C8Z0ChX5tkk0ULsWk4Qc5yUyWhYZkIaAFTMQFoaIbr8FVPylYJfrDL5q7q1eBAKDAqa
hNHxFVbhoYzmw83BybxENiuuu6Ci6xwmJoyUWSLa3F5FE8sr70ZphxW/3THc6+OOEgphhpUNvvQ9
Xrux5psg+1FpKrQ8+qJ6vb/CL5dxpYtqUYLWNLUS41DrXoxE7TkbeKlmy8/OJLqXH3usQANWfAcw
vG+a3F2+H28ZDu6VgPb9WIXLMGUvD3LifFlGXFM4owJfgfmhgk6PdtK9PUYMS24IrBSpaxqbrLzd
DFLeTUmKP3BSjUWdtr49XnOz/1SDyiTUk03CRZNk/WBCnReXbTd4lHcxK9fFx0NXi/8MNSsU2dw4
zPpsxr3o4oo9sKy9dkRFHX6oPdoS8K88ZHo2MGQKvkYLK1ntsN2FEWZl81+pJs/fmdhwg/OAdD0S
Q0qvFqwlUvRRT3YCacl+ZwSGf3dpYvWsuK1FL47Scm5lOX2XH2QKlrRi0jOQGKNhSbiuKTlAmNzK
WXF8fbBZoRFaRYXHdSpD1BnWZ79h0Ts7ngivmVJ5cIt8B5g3HQ4bTZOxjGFyEa9BzXc8UPLc5pdS
mVHaFatffrgFx0Zdkj6VwPAgnU0FSyw2j/0y42PVMCjhjHME1Eia3jIA0R/It8syHkL441dZyBO7
2kkJLcxs2R1kJo5mZI+XNFa9Pabga+xpMfEOdJK9hr3qgEsP8P2gvOZMIvhmbbn5NdPN1o+bcn41
2W9G/ygv2X471ijZzuEE2KNfHrCZsNURUO51Q8uHvuNk2/JeRDIM1YR/VcRz/a5IsB5qksLKG7EA
B88BZZuZfS3UI3Ykyg14sYDtOzNAs6zAxSwApUXWZcyneRjC8wkqtBPqfqcp5+S6erBc08oM//1j
jO06Jsu22PEiriXix7XmIZ4GEw85JZEZK4B9rpDVHshVyEXXls/1V9ZNfvj8V/+pFTdNV0btUaHG
m0J2fzeTgO38+dCl2wKNtjRNo5JHt5opUq8re6OeMLv3+0YzdI5JRjaSssaKs1LxGqDpEYqiBubD
vzVnyoWvVa7uCHNVLsjQp4GEU65UhlFgjA3BcE1NBNfi2yQGPgeXYao3yDHaL1NE/7TiWlT/H3M4
7Js18zK3QfyqdhuQRsYpNHG2PIp1R68hN4Tc4RjOTXan/5rbMpdRF2V4pOdWFupIkoIathFxHYsx
lOr/YpXbnfID21ZxHvmm6xP11z2zH7StvOwPzgp8JXNdtjO3j7+Wgr3QHdjt6ns07FMcj8ZA22XF
Tc9QINd8+FF/o4kQkbnM+3SzxOp5HkX459yw8UNWx/WiplR+DubUnvrXzpeie90hfNOn0+QB81MN
DxGffLPw3OSiVRauymE7aYt0eQjUkSGkpHrX5Vzv35xGvJrmM5ep+vcd4x8Dy5ZjDuimK4NND+iA
Wn82/e7JyeUPaeuaY/eq+RGDapFtGt1WR2xzJKAO3TpbyvzHWjC55FjRkUsNvHd8AqEl2MpkODnq
gIrHMlpgOoz7j+UflUEklkdk+eEfG1FbQAzMsSLxWmDxq6ouwQB5Ul26HC9+jBcVhZUofPVALPtX
8S4AK5d+2IPP3oWgq4UivFlqxdeULtLcsSNuw1svGood5mUsJUnAbQgvc+cAqW6VA2DhF2Zd3xIL
j4M8gyi9NyddZcrinWV+Wn8cgLmSFWBcyZp+cqiWSM4TyJAtTQ2xzsmryfCEWW0RK96TerYiFEyR
lAsHFou54nfaYOzV0pKsdSAUrpmgU0SaqM0Ic2wz4MUVW/m3op6vWsZOlQ9dVpKvCBS4uBCJXoYR
Ws+fUGt/d//KGIlZ0HaVyqMX41Le7AbOPZoELSVFySO++qJiiholbLVm3xjYXxw9cuGtIGdq5HBP
XkNh1UKNEj16DPlyavoTazQmBXe1XmcZlXbIDWIb4zfkrIv59jaaAyD/+WSEbnp0FYsNVZ2HtZVk
Y0h0PXah3RWjsAqNapgrf2X0rgSkvPfFtXKx6v22R/AHE9/ncAX7eb7VS+6LzK/RSvUMWouNCiyJ
A96K60Hqwt0uH3GhS60isULMpYV8clMKdDwHqaAbZpm2zVHo9NVkQWEpf6Ovu1thWv08Z2h6FTCd
WzokFBgShTy3eNJ7XMnEJw3+8/V8XzWGcpChI+zIpMrxr2jR8T9U6AC1ccuQ59xTaEAxRpHd5rgs
P5Md3ZAWEXwsuu9a7mSxPjFQ7lQdvZF/cM6uOUpeZJwqaLA37rKiw6mHldokzTU8drOtSayHjUQQ
58vPt09b10OxK9dNzwmpCxKoLpJmruwHm5ldUdnhpW9gbChnLHj/0AGW/8s1mwsvSROLuZH+OMU3
hR9aFzvoXs0N3HWlvhw1RbtKwZ2HjRqp8EheMfVpUG0trRlOk/Zmxerod1axRsP7/CZ+a1nwvimV
gWgeU9Xsnz9Pl6gyckyWXzB/qJVoqE8X3q434BGsWLtyl8KH38UAgF0YHWtZqSgcEsmLzpUFUGaj
m/dgK/SFuSmmJpRvbUXYCtQ+5ITVHecz8bU/OCKSVfyPsGn+2ZWURxc9fUhgceCRPPq6eQU7BZdO
HBFpoqAeBsIEG+jsH3qzP7yJrF2YZItYljXqflP/CNQPg86iKJHbGZWbQ+JAfUiYzutdHzumV3/g
rZh5bEpMs/ATC6A7kn/gpZg+PxWf1u5aG2sLd/f2uNV4kvn8Ck1Uo4h448r2wkzP1FLdUA4WEPB+
7kw8BVhQF2qSxTZVo/G8fBtPnw9TYA/kSdgXZGrcdv0KZ2hSmH9rJe6oZXXoRJtAdn+UkFFfZshA
olzgPV1ZV82jfFFdLdu1dis21CXqRaIb80EVzYEuRGZG/REo/nhejVd1d0goOH+znTb3hjddTQDR
2+aHUXCD4uDK/qMxTxEDU6jC7IXmzmY2/9erCFmHPGHm/M/TaQkk9uxgX2sspb4FLP94CPZZTq1R
8lWLFBweNs3ppUg+5ibZ5fLxE1Qtg3uqxpdJUTH6h479M2IPPQyUc42ierZFLKNLd+j3Xf7eIAhp
V4TFw87LiiqXURCxnExvrxUQNAui5FxWHVv1PJk2RXJxuvuZ/DAwRnmNuWbXaVS8b43LjjpX3t83
cH92DOI1wSAIXIdaf2tA0uAl75cQxl5K8lwM1jyQOTfYPa4BGkM+qwhTWc+NaOKq4ZyJX++Xk4cz
eMFu/Nq/e31jCdKGuyYk1znFDLcZQUqfTXZVMyuBrsnDZS4/sld62sUUsV4whdn0VKcPFONntmnV
qQfmSt0UpqGSMrSYkqVTKRq2wRvkhxe8mO84ZjM5Kjc7u+I4zAkST1l0F/lP7IIR9lMW7Sa13sAy
4ZjvOkMQciFY4oMT+cN1I6fK5NdpiWf8lXwZYCVZrD6a5N4Ftydqc/RHADMnsmRMTMZK16/e5S2m
DNlAP8CBwsuBB1fTvSYsnZBmf2dST49Cu7qxh21+cSyM7P7iExd4kfVNRvwhczpy5iIHqSPLyOfQ
Q9zPrmHD6z/x7ci2CRJD5hkjmDjpZ0bprbnMqS2xsZ0RbU+roZCZ0YYIa+TbBR6ydQrL373tzh91
3rw6Bz27U6kAOckP6F7dP9mR/QSdHVyqWvGrjGrIFg06+uIxLA55IBwgJd4Qt3Vl31Ti0JDJbxjM
5EcGDoPKFqz/4mclsPW/n/Ia49kLNErlc0YGZMPLdTXiS+1Rkr9d+I5jUhKLszzKDaWmM8vybF4W
DJ+Pbhtm59gRRqvoqeAZ0stxRsTulV6HifKTnxuZZtGvzjB9dYabDz0ae+eAhR10dfgYaM5b65SK
OTbaJwxKS2Jp2sUdBPBhD/CEnxJX6j3kGHDo6bsrvdy8JsotGQ1FlcqSwrk/r2rkxA9Lmsa1KWCs
Ttryi/XLWrHVzlS5UiHqrgAi01TDus1RnbpoPqaLRDX+J84LAWtOcNtZrQH1SHwklgN0VKir1GYK
8ZHGnhClB+7kZHwHRnHoqk6JoAuFJTZ/WMGbRZpgFEb6D1cPpZCluM0KQvyU/tWB5XgsoeLs6r6H
cSzOXdltY6Sl8H8X+BbPP9+4z2xE1ktU7LEGnFjmKiku98wz5ua96ZyN1XIMQ9RHNx2oH+XuWp+N
pQnPLWOd8bnkDAD4rOhGCQgtV2EN+DTpbsMs5QtMxxlKbHWHk0QRaPPJAaXelJGCZgFGiiVcH6xV
V9EyOAtfPOJtFvZIxnRHPfRQeyOSOCLX6l6BgJQHTW4I/t0OP0ZvSlsQalziOTPKGaCTtY9bwLkB
EYOe08+iyp/yZ7C0jIrxzHxrpyEh2CnwxYFC7qlkzXOYZzNcKuGRND/mcHQrT7XXnMbH3Z/c1Bc/
EMcpozzvTpd5dCyCQFgPasJfzIzG/gAhiPd3INTJg6UieZYpcTtLFhCg4QPpZvDJD/IEgl/QX5Mn
0akjtkk/HzTyM9SCQEZ0HJOQriplpBPjBcJx+o2Y1c3shnYY2pc0LzGtndQXdmd5qqUlMlQ5mRPi
jbJzQy20ZQjmYmG64TqI3g7qcRV64OgBSWTrtd9oM3CD9pXfDgxk+sTN+K9PsnuC9UwfcuN+2y/e
tpl61FRoMiq7PYzUClowjBOjQ9VKGchJFTHPR41RhGJaKvvXC+2yQrZAc2tX7wKXewOsw6Qq3uHl
BVO7Z0DSkwswwdWcroc9Lqu6cDNukEPmFB2TEpF0vYTWKseD4l7gEJoMcPIdgflpj5/rUryCt1ZG
HITLEqOPRlbRsR90so7T04vRSg7T9lu0RpPj5Kek3igEXzkvYr30jntd7yZFT5vPJNMUOSkEZJma
/r23Z8Zu5JCnLsqYv6/Jp3WOdVH/7v0W54mUwcppAlPZAE0MKHcWuHkh55WAZbczVnSo1KOAYmhI
qhb6NjMINBJF5nQoRWwFNUp2LlN9zgUtltrHGc8BK6FaBtpxatJM61XML7gbEN+yZ+4iL9mFiRR6
ind/DWGkHhdWqMfF5SnVn7UWGEUAMMlBihdXvedtWlnfuTUB97IufSIvamgJwQIVbjhEtNdl4VhC
iBPiT5aP7hZOf0T/bCyBxHajW/FN+oI4lhSmnhbHqVtMg3638Y1bC1Yd9TA73YwVLV+2nVPC2UDI
a7iCJhzJ7TEcRZ7f2AtvZwQV1Tu4fcGQF/aVPae3KS5JqOBthIIsdBvSYTaVkDOs7SYrMf7eaDqs
tFXK+YREljU9/9i/bvwsM2DY5geOhrIbqq8Z/xRC+Jjrf3MTQ2r3nkNTBPhEoE29uhnjDRnUYT2g
epP8WuwTqvXFK2ov60i0kJMYSBozsUglzBIdrgj1alntnC86oubfaccyV5vqxvP9snCjCwuP8PgZ
MmgyH29RX3IwZDQuUnWT0lik+t3NC8lWx9dy5IPS9iyBfJBxpSSVl4+9JEEVVBm52ACRL+krdBrO
EbE1ecdgBsFFUHyPYWRzaMIoaxiDP1jG4GimYKegT3tcfrw1y93SdmelPzl3E6SGEacm5frxmv6A
haoLq6CMKQKHTdj1RmaM75yxR468b4DnbDwdSUvo1TfZUY+dPy+yLjzrzMnxbalE2fXUzJc4Q+Yp
tzhLavVU9IzAlEU/71iJxmpLluGmWjNYqtz3q9L70kxNDgr1/v1tzQtjZ4+0kht/hiEAGsv5yGJj
9+SIV1l2h2OYrpEhOcN6SDgjjWrrSeqQPVTM6nnktV8P6VvmCyPnS0LTmajk8LbFqRnrrfJsA8Sh
4Ad6VL4qjs0KuRLJdWbtXb6OLXI/OGEYGc5yK0oYvxP1V/lospO4wdtHfrnTdRKcZoMcYGbBWEsG
SGd2kjXZGvNBqOe6GV6N6saoM4hwiGt6D4CzkzpiJwXz7ar5J2/Rew0DhJzpDSTv8yMB7Lom880x
9kN44QZxonZgL+qTYWUfIlE/kA8qySmrVlEDU6bNpCC/mWbKjMVb94utR1dirxK3KeP99lefTl8Y
hHF1Vm3Pxtb8VqSjH8ZV16zblH+CKbQcFYnEaZoUXOjIctCiFSiWaruG9T9LbY5PNtaG9P6gmuzs
bdyb94TvlztWbFtTKqDklqh402KH5g2pRI0ly5XEPJNLwM6oApM9mgOlO1OFGWp8YClKYkLFRJ3a
yT9axB3fUp0qcCoCVHVYlxzeg6hCF6AfDFy7Hg/hZ4q0OAGhzhmNrHUwtE5PnbqKacBB3mP81Y2g
CP6rchfj5M2m9Ky0yt4tIXNv0ltMTmyqvkG4ubFyZkgzOnazIqc3tKFqVLnuLybsPbgOSR1e9/zg
Gkq8S0brjSd7Q5UZPnJAtZgJ2cVkn5CX3e6N/wY5sZw6NDswHETn8rUt1XZMeM+roAtibIhpWnmG
UTCQVGnuSLed1mRArmq3oVS2WNickBIKaBmkthaIw3D95QYEUobEX5BLsTvGTUvdfQPsOxnMZABr
nvb0Vohk+06T7W5FEfiv9DTSGFYQMf0iNuijjpM10y/Bo7nlT3sigEHPTIbqyuuwt2Rw88/Qm5AR
5GgmCgY2yp20CAKSgtyD+iR1wthNkYjWOnawbcsfZyD/uj4FB92ueXJ1T55zqwUzlP/2ZdzZHdJw
cbE2JXq1OZM3MygoQpy2cDcNLkYBoMQ59gDj3FkurRbXzZiw51E8D6L1DHrZ1W/Z2VpoxwXVniqJ
rLI4H6poBWtCnyCUsa/brzVeKWKOHbwnLLNZjqchmIeqoIGP2SqBDwCtXsIOfFRCjd94pkL/ldYW
Dq864Ssau9NzW0PomtkAPyEPd9WxsOm9hnXDQMFD+og9pFwruZCcY/RZNfd4YNEqBeW7kjjMf9+q
MNK8a4OOSKDKZk/X1B/sNGI3qi5OoVqaTjdLWcvKpCq0+HlXpNLvzWvYje9Uy0jO9wpD4lk+2XSI
1IPp2eUb+raDHcoW4fg5hllrBTDgzdA2fZSyc0scTP01fFLsUok0CsQ3paQIygBJXWmDi2BBqfqI
We9Q+TVamzOdVxhbcVWk0sDpBwCjhMIb4L8rlbUQo4Hu0SqHcqeYkgUwqjdLG1A6azzjAa9mz9/d
XHuanULzGrF02xZ+dR/i+qkyTnqYPDLnBgzFo4SCqdAIv91fmXXHdyHgQSWQDjHBk2d4Ia4lCJqE
KO+juOY7pXf/yFvlrPTOo/1qmtMinpH3zbITHSVLL0V/NrhuGUnP8XFWELtp5hMLpm84ZsBDrU8+
4pHJy89z6Dsi0EwtRd41XPfFmQbbiA0F0CTLAp7aAIJc0IbH5VZrNbRY7lmnzduBZNOiqXbx85cn
Z37aciDX3Su/uT6F5BCajK5LJ1wlN+umGi4aJFuZ8wthymrAFuEM4S5OUTB45kCERsm1/oO0abv7
mb3mGkdTINmhgTxgkzZnLudpV6XHw32Qr2nQGdnYDFMhX6e6x0OuQ5pcUmk8n+TglOwrYsSBN+H6
pESLVZotrFj8daitrXCMwJRgw8yh6Hzne798dAGJ68J8SQHT5H4vuzP3J1l3NXzqtcnc1ap1E7XY
B5LRJpgJBmbtqvNI7q7iOVIfN/KNHkMlKdFjnI5twwkXbO36RSQbs2i/4RB5kkpAtPXhUcBMcMAC
hrRhVPenoe4p3TKMzcK5B4vJz8LzIIOWu/VrsIuJh3Ufl0BWsSZ2FUi67Pr4ipp9nKIjzk/mND0+
RTaIuemBWyq7d+HTIrOYPRXEkabKSifvJBXqgLwbbnFR/DLOXmxo1+IWjvL63TZ2PMPjHf7x1L0n
z6eCjUOKbYFTEf/bvv7k0i7g0iz88LI7uw9fk2/Unsb7zi8dlEA80wImn4c9PJg6JjRo7g2HVgy4
AsPuge1D2QrADCGArr5EhtAPpAhVyGru1PMzew0CqK1d7owChIzLVeas6+i7jF1MuSvTgVaToekn
Wpj60/WKbjxwen18pPlpe2tF5JsRpQqZZ8LhjPmrQnqiQrNqqZp0pOBZFmTP4ZNvM7zpHbeH2kDt
j2y23xo9CqQI3CeEJlZBqXgZYYq96EAW16JwuCAHkU8MqHw47b+0NsymGpa+f9RtpvYKkSfeMrce
r7bZhXVaZFhYbtyn1XAIWz5DJIqHlm4zrJ0rRU7F6cOJC3opnMDvpVqxdjniFgMGBl9Pb+uJG24c
adKd3/wkPQmq84ZjqI5UtggHGzjCUjdtSuTqLJHAOxy5RvU7MqvGBi8CR5NLAadoAghImiy484T+
j+ueqHPOVcgALIIrVmjQiksmd+3LOowwX44NMp4+40NM6VsptROjKeS5D+5hAY5RORtaWfd/SU9c
yhS5A0bX1PiFCzhsXH+yNZbSZ1oN/v9EOAs8+zxGg15hdGoo33b6+68MenvjxTYAI08UfjVq62fI
SKqdgyDNr7EiO6AbQ2DZKzmCcC3Qo2r+U6RLLCLIAiUYoQ6evxymSW6tPHoPwA63vK0EMGDBHhT6
fT8skYOGGgJFn8aaW2eANMMJ3wZXiLeQCCIruFY080nUAoFxm0nHyb4ZupMZLn/74WmVIQ13kbPG
fme6PZS4MYER79EjIsDcxAVsijg1IcgwJCp20Yn7MwxNlEG1pSUWSgClp95m+CJQEEH2UbUSYCWz
zKDsR5A9oLtbHgcMRm611lR+U/11HqzkpBNUks8zzehHAnp3DmALMZXwimqnq3Xqg1IZrkymleWI
tvEQmZzbmZUlcoDs17TWNjueQV65pHELtfvKpQY4araBC31zvYbSx34VP0SBnh2jak+emUn8/nt3
flJyG/JtbXJjGk/jAK17d8bZi+FPsPZALfK1u677t/3bruWhJOcUXG7nroQRf6+DFgFjbY1Fu+aC
PsHRWaqJHo7hin6VgCBweJFHijMsVHKKy5Pcch/qk8o8/p9gBGZeJxnwyh9tGOxvKU/xCieTOG/h
CVmkbiaMgEfJc7h5PvdSyoye/18EnN23kuSsXgjSYjD7+ii/kAFLla7e0vq+7uYGStnH7b9l8/yp
zo+biqdNOmMjG14Tr1i+z1TRAnCX00w+dPj2pl5A88y1rYPuWoXYH5nhoLv5xdG9F4pPQHbuwgiK
LfqD7aszANU6polNJPUw0JUbkb8k7mBmUt6GnFGEPlnTOzlBJuTcq6GcWRe7hAJkrY2f7FR+SlL+
e0m5CerV94JUtCl8uEGT7RG8Fszhvf+qFxzuILyLiDYmtLvANPtzuWiullzGP4aGWPeR6n3WyLKB
2zC0R49C4CAP3b3OiMMdYRUamKRAWtULYPOxZDwqTC+SHUQOhegDqQArOx5fxEnbQRVuc8Ys3jLh
RTJbR2k7EmkvKpmuJiu9KPP17BB+XGXL9LwMx6ka8uhrZTxQCVCiZ+5UEAuhwQTrdNfmj3x7HwX4
H/zz7YfVFDUVjt6wWVGlmYvQh0s9WpjG6E4056gGKRrVVnuNs7rpTbWeCAxoy29UavtlJYX9wH2h
yvBfCdt44qb7iZJ9C9/mk2HZ4tOxDG/O+TMmzlX7slVKXerXKRAAw06b5bytpkD4Mtwt2o7IMDAg
6RMAw0zrdJOb9iR0tET2HC30a+OTaXVr4x8CuIkjrBCUDgMEGDRBE1mobq1q6kkR03QqHCNrcdHq
QBxBsurU1wPWq7aIVj/zuXyJByZgjnFwyteyZMzlU0TfhRpoT99ZaDqknJ2LUI3V2ZQfKnGoJ12h
u/+W+EqxKAvu39JPzKkdAyMSCdG1GkDskVv4hkag0EyKuXJgXFqKfvWdCZap8daWj/hK1B5uiPUq
B1pMVmvzCQOECRZlseC8a+hMmVujkN/bzB7PvYb7NzGUWgrodcd6UKLU9MnaO0W2SJ4pzxoqsECy
MbePhJopsxBvKFL9Md7avwCZcLJqEIJKFR7U+SuMZjBB+N6M0qMCmMeCiv719kEsK2Y9SgBlnus4
pW1fL1dwayEO9g6edA5FTXY47BvD7xh1aLduA2kjcb7O83MW1/9QhjpHkFfFuwF7FeybUkv9wlQ4
7o3ln/3hLzQf+JZR/xINP7h/eaadOmX6zPMv4H9UEnIx+ImQ1LxvPSdcoq+MR7mOP8Ir3/ACFgqx
kvEgcJlIytnju4mgPORKdtyKaKGuEB4XMiCQLotD6E45XM/bDgPwUUOzJwcQzJLEhemiGt/O5iuq
YD0cHSkbNsZ9+qtpYbbbeIvNpxJNulWi4Skn5UgQM9LUsaREsFSjHGBQii/LZAPtsxpK23Q2PwBC
EjMC7c5rCl5K89CQ1/6UbFh+k5BH1cXJ1hHuAP9JvA0a7PBCxx6pAllv7bdkHwVMtC+N2Qdya5Pj
gAJQg/AMcuncf3zK/sZWkm5/WV18dbpAN0OVUstNNyPj/5OosSeCg8o5H4kyi+Gj5SGcnlQFcTYd
1qEc7O/Kt5wFi7PQ7lJoTTZlaARp6tGme/+ACtGejY6J483hfIau9NibZ1KmuTas4kIA5zU66HJ6
o+coPopHO/qhCiFnWHwJbSq5Wxi+5ZbzY3ZuOu6WJshuGvVSr6J76O9x1kGb/komv1QB0xRWc9ZX
X8NC1bntLJ9bIzraYg8HNABY0Kzgh+Gf93//H58yjWia9zOAqFEKY0jQrvIyF7F3Ogu7VIeu8GMy
UPCrx706JQDILFy0OPrK7zy+GKu0/GzM7Du7xtWOgKfQleX/3u2OHi8Uu6bD266lIyWlT+kiqI14
OKVGIUkXWEprg/eUe9UIh46JUa2000JBlnoeHcO9m7tDdJ+eBjyajLA01tmU9MrDIg8FNbpdklKs
Aqw1B9V33t77MsvKmMNgNbubHKiJY1qlo5vxC6lIry6ewERKfWzorOqoywcj2nEss5QmdYPodBKk
3Pjv/oRR2hxnNeOFm8VgjcwNJlfrkdKgrbb9ZdwYBC1sVSQv0G7BNDRuRWDl4VWECIhhomukR6zn
c4T5laCAh1yC5FxNXThFyd4zPzkOTRFcU9eFhP309zp/qLUhHf1em3CR2273eXUAHcRuwHFInOJL
h7zEVCGxV4uyVDhDgM4epm6crwCN8mmrNGjGJcT88bbTcfcVoXOHPP0rbHB1TjxHIYiJ4e3u+ozf
F5ev4j7UJEVW2biBs7FcEFrZt/eK3cHul4T0AHYPcT5fEv/vdIpQJnsU3AMoYoZH1Ef9dqsIRN6I
wvlZefBcb8zp4oq6wnsB5ytwzKzEq0rl76cfWn0nRoM5IIWi3a+7bWAzJaFX5s2RLqmwdcpiPiF0
DT2PQIFw5ZXANGML5SOZthx1Bvy9oL7+HyqlA/0daoftkLQsscvQiwUKeUA840A+1tkPGFqhKe9t
Ofu0mf2m97UvJQAPR0w91cy0XNxY36tWDBjBPilXWmln25U7xfSjNEeH5XG92GzzJ74n9avkDYvj
Rf4vzXqnYBVFuEwdeZ3WVQ6LmGYxrKujjck6izE03zoUugCpf2N7XUudhwZPV4hte3o9X8ESSkn1
t0UCM+DQZnqgbdmrIw6jeyyD98s+c0JztpEgu6Ifx8ekLFilgj5cm7K9rBK6MvoySmsvRo4/EaQT
ejd7kpX3b4WfVjfnhbinn73pIjgH9YG5fowgT4sGuEL0eH+ByRO+u6n4P71Uc8j4o5/KPpaKlANs
3IeAFN0WdLQlMTurNmLmUXEg9nCiFwW73+1OaQOhuWXA1e+L3drRhBe+N1ee5GrES48GNacTPznk
MQgexZMYv8fLmtpZliBOlPc6fwBEuJ44yq2/1mqwMXJTmfLRCDqeSlOFJZkP9MPLznXsxTtBD4EW
tavqsNQTLCx7T+uwCo1ecHDM4Gci/cmtNC/x+2z5PALsXF4i+KHE9Rch72XZ7oPmg4ocfRkWX+E7
0ef94MCXpuZemN5Zi+K5pTWL7g/xz93gQfyNtVhCNjPRkRmLR/d5VPKoI9m2lzBoDM6cEnhlQNT6
b5bY+iB0zVUOVj5vuwsjp6Ubf1gAFz03Vj1z8h4gtByBBycxThxX1mhkpk+uQDLOwSKuWbkqax+/
yKX3Vgb6b8HPxuZNODWL+v4ikjZijn2Nk+urYM5TS9Ji0yDkXHam8eAh7RbpCfx8GI8x4dKzuNg+
gYIPwET0Itl5FldLhgwhNs5UbteYK80Uq6YISAYtGp8VWQrXD8KEophheDTR6YYswoXgkdPz0WYU
MtRBVcsBOyiahhn643roJow3Qam60RIOTr69GJbyRreAOGY6Eaqy7iBn2/L4q2Qdya1eQcDFxxBL
A2e2uudRVdrNNUqPl9wJKgfAViI9+keDSIg7/51ppITZYto7dbAMhJoSKUCmNm+xgclUJaZfwxrj
iSuvEOIcFz5RcvutVQgokvUm6e7+HKPqJ9Ra2nyfC2z0yGmEULLZS6a5p4PIuz0aSeQpvhtHu2p4
px7HsbLFDj3IFy6IMY/wDKDhoehLx38/3F6xhfo4SFRtwQyugUcRaSXKyE2Ne9VF5emX5xLoK+Nv
eZhqkR69ACxgcW8VmOibW/c2XiXGHscxKmkRydXS1i1LL3GjPCFEHxBtswjRSSyDgcRfZzciCKo5
DsJNPzgUMBjp27aA5uzZ3KLsUi66DacO0BYvy0K7dcS0p8Ddz9PKjUqtZTbC2xVQvWD8cG3YsPrc
BTn5vftWJV3FCnK5H5DetWn1ED6XvX/8uGzXn97hMsPYtdXPioEOXqY7TRJb5G2BZBZtcfHDtfLN
QD80MvRccRdPBk07TfNWH5ZgvDMIFsAtQGVvQcckazLiL+kU+/j0rlqP+tHTMQFLWoTx07kWPKDz
fnndBhViXyktJNAxuZ2zAqiTQKqrVTGxYX+BUDGjIZUT2FcqjhfN0G4WWF1h8lCCLN4i3ugfnNO7
z2ihqg1AJksQfDVyzu/0NQUTtRN9Y0ad/ry5+qgIcy5s6Ldje/8IAtWai9+q7mpojvgjkYmkEydK
HNYT1xFOpw+LyFywm1Hx6EkGPVusZ4gjUS3+51Du2y5D/aiZtbRo0Vnb+GdS+AW1TfG4NYAaTfrx
qj3uFUl7OhWPHSnrh7PVwtbeXr0cwQPslZvUeZgW1WQCd3lWddiKz7srFBE/wf8CnwN1AU2pMMQX
ipOLoXY3b+qiOnJqyHVAlv/+F9PGrMdityl5sl7rt9Sg69Q911vBH4AlrcdUvkr5OBBxki+cmP1x
BDtqk0sDn/jqCdGs0Vz0t0PApUfeAH1jQawQWuS5L4ULQGLB4gxWJ194rI3drlrD7SSRgaDuix/x
TpOruI1I8qkw6p+bd/DUrv8XCaUGFaKhqVVCEpSsbCHfABbj7wvw0Xu11iU76hFzid0nVLc5oxrO
32eAdmPBFuX++9mJfPrIJmzhSFfUmx+y4SAk6cD0ypnMxzxO3efxpu+GTC/wNjok4HZsz8De0Wpe
86tIbebhi9Fo2WBwNvHxgywvmllQU2AQKZ+SZ7nLRJeB3UwuiR5xJGi2peA2n3Ed9T5ba2r3vivz
yIc7cBUh0xWu6IHXlFYaIGJ8fZ0gtoqhKWjJ38dl5nznYxFP5Y7Z+DCrRiPQmB0C0gusYCALlaQn
Ts5nEIly/wBdA14j+HdcGoorzUAbdS0oXf2Q8oqmj5UyTHtmR17oxApX3glJxgvq1Y5CFExE7G8o
Hy40AOr9ncInh52loP+Yone4ol/qkuG5XIrYXVGytmPBpJN50NFuj7fxkFbi6nN8+ueyB1KHRHbT
nYvjuKBQU2/uDTEtke7Kl79dlN3T8Rv8EldlAiMvYEKEfmePHsmnIpJQW+ur5olqEWohb+Spqn0c
A6u++2uTUSKzW2e175JylJS1B55l+chdlXkTv2SqvE3XYq6dwTG2C1uTN4GHv+mFFKg+2O5oJDks
5YgamK6mFIy31T1s605oEQ1nmbToGNv4vQjUaaYX6f5kxuOD1K8R5mkwVixusQhjAR7j0xdAPBMy
Vg7e4e9YidB826O9vzS/1hib/r+avCuPEP+7lagcy0JKwg3SX2x+oOM6l3MLUpU21h+K+J/sy32B
YcJVKvTAgkApj9/XxK6YUr8VGmgSuvf89JQA56mqD6ArZtco6ZlkTU3D7Vm5ItEaDs5I4izlbloU
SKdgzkQ0heJqcjIb6HNK2FGJC/hT3Lns2iIgyDqU3slZBZrODqnLymI+4fmAyOQKSJQ1ablTuWYE
sXTaey3QrVNTdQ2AJNLncY55qNTSwM/aVjNPttQs22LgmRjy8aX+dTsRL7YCWPToV1CHaGTIb2qC
f5+3KmWKX5vnJZXJT3yq6tQ13ZDNr/kXkIwY7ZhGnmmD/OKi+xgyQogzGLlE6B2Pnq+yFlKzG6BQ
/H7z31wzrD1ewJu8GekvxOpsDU8XoXLkP25GAWClgw4fVsjMNYJEYwelO5cZ9If7iDamWh6vvFlh
zneok31ZULUIjpo/zMxBUGM7PFDCVAyJ9yDnzWrZfROHM86cK/cnnwCnGP0QCD6r1EORQxGC3CeB
UoymferpmQ06WOZi7ysnpgbFswmmk4BXMZW+Ze+NZZ2lHuO1EDfhiNIk2To/cLxz3Xg5F1SkZ0cO
cC6UPaHnT4PWVTifVkHZFCECRD14IJrqe1JNMS0Za/z2bD6eJKwnNN+z75UJjSgpHO0C0UIO7xga
8ouUQ1j4wQf7zzmECj4MsCd0utn6LfaFzNuhBBnSzZ+TAlqpO9gOWA3WnJzQmN2sy4ZbEjHM527D
GWDA9X7keo8gMnGuge+WxVUGzPrrczRQdvOjBXGUyB2qs2Me5Gbu/g/+FQujzbQfe33Prlr8+m0l
2CKu032sQnSmitdISNBu3rHBYDrz5sdvMunsRWDW0k833VmMFg1JrdE8M9nvfLHJv6J9Mvin2xEp
laZjebqu6Gu2+k5jh0NwCIuDfu9bOAduPoXemjT8hw4e/QUk7oEVfGzYMCbr0/UXzTqF7GqnNzTj
O+WvZfp6e9kGV7lvHJwFY6VR8V+TeTmMO8q4zSGA16FS96P7m6DEfoMCDCZbneKPMdrX/X4Xks4v
huMWAxKdhdjqblpoLtRJ5ngmLxa8/YssNGImqL/n5IsQHdCLQoRkifQ8DrgHPYE8Of1Q5Tqf+j+t
dQLwq8v0rBqiZoD+ch1tyyBldXVJaplfPLmix/SsIWDTItI9LOIXmUnVhY+4Wk42hOVp3AAVNs0e
EzLXXJSvOc9vnvHJI8H3mj4mUKILYKmHqn/uAdirIP0x5ttaLiEEBZncH3dMhhLpDyGcs+EroB+P
w1j02HcR9k8EmtidnqMsBZphsD8bYbpmIDihrQh4FvPIXRDTRFl++d4BzGQ2aXHI65K9eWZDrqGP
DrNGzyPLWm6yBh2LeifKezjQvjjtW//X6/sRm/Kti3c36Z75/1gXPi+ZcBUv3qtATCgRDs5kLmEm
5wdb9a+40jO4/oDu+EqK9vGfAG9DM9/KI99ZR3TKMm9F/HUXQy/ro670rDo8llOYUACq274F2Kwq
HxRnyRpxkGsDY248dE4djAmHCOGbw6aBSAq2+0BMsDq9hm3KsziTHOMoLV4RbyhtCAK4edBHu4Du
AwjyzO02dgikxognkTOFqggPwkrhurcO4vofODn8HVMh63qoFIQmmrH4wNY/fgFyUNvxwaJUaGxv
8eGXOXYJuDAcKf+/J0qbEaA2rBzfuxsnRszM0rWwuM2WtT4QzcS520RF2zJhUQHk5/oWz//vyGhF
0mRoaDBsTGmZLyPQZBXBuq0XodOSFrusWjc/j/GPJBWn0ha/3JmHw8Pc4sWpkjICfRm9A8yOqmiH
h+HjNL4AmG6LiInmzLk2qZcngis5IgdIpcyRWhX0OYv+fDK4TAqrGoGxc2yl/8+AxBjxAhHzrYVE
d7ffCZ7QsRKuXlRYpNuOR89gF3N4b2OMbiHlMtVau4rRE3Vy4S9toJuAz9zaEAxyXLjEpa2+U4z3
WY3eMi9nGj//yElu2UB6jlbAMbEHhe++PUM1J7bbA3X0HRk4Kq5lMy3FfqvKu2VFaiM237maIxc/
S5gLm8rhntm2miYL8JUeH7cjDb/i0Kfqb1MUV/u6l/ja/flG3TFvcZkEOROXgz4Uw/P/KiBjHxTq
st472kRwz15s7fRuWuaFfQVa32108Sy9f24LRcEwbq/mBbgNamYMRTQpNeuzg79NGsfLJC7RI4k9
/0whw506B81mfwo3TKsAo4kOGYess1nERC9O+UEuaJR+qVOjfPK5/FU2FVoAR8TUVX9JRLDGwNPR
SREo1vA+nXfBKueE99wMIafFsZ+lKSS51/1ebMjDYxAlhlvNbGdewMFASGbSv7LqFbpVM1rRBFr+
/5rPyoVRdcq45mx6dxTsgnHGwOcsNskdtXq4hdI6DNYs2m0LZzRyeAaBX/QFpaGA/eA5iCv5qDsJ
6hcElAq6Zjl/QQv4CS6K6M+hv2fqN3YlKbLlWnKvXHwPEy/WET1/P8oe2O0JYFD0mw4GcmM7SYU+
++QxF9KM8EUzyWvhHBrAFf/RPY+Hjhtf/sz+vg1eoEhizUdaGF79Kc19xFctvBQGV60lgFQjkLuG
BtwqSbGCvYYj/uJzzDuV2NB/EWj5hKd1JiVh86icC60NeX3NeH2Bvmb2UtvzPdwrN+UCkifLG9sK
4l4Dcj0HdIO7gTHCulkbKzmtOQsVdIEBMSFw6NW1xlaXcEyoPGC2Koa3WBDL1ICqco7tgz8jhXgd
VfTwybuKdwpAETcRJ5Xhn1lcgGxOYrgXox4RtuDZsGZbiocFaebHchv5kI3Ugk0DzN8OeYq00X15
zXxVxs+Ly+OBWNoGHp8W3X0Ii8fT5QrfXINSrSEfbIO3BM5GSXTCJ43AX+TXjV/yD9Zhf7Njk9hI
cjz+gRokDP1G8Td0IDRQ5lydi4zb5pOn8zIq2BYJmCad72dJuOe32q2ZOhLp34UL/S0Ky5fq461m
XJu+JT6Kaig48+OsqhKdvozLU6ii6W2a4EFBvOyaSx9IMVINm3lABJ9NoOCSt/mQE6Br//V1BT9T
/fS7a+EUu2bISXBrYUqcK5YJqDmyZi5pm8k9VETroKRn4AuAQDdwrll1DY6ibY/Bv+SdQVEdftA3
dwGwDlLRmH+NX8TG2b+QhF6aGcoo6e/ckgyZzoUhaGNhbyGiajQJZoMg/RN5AC/ZNw+oqXGLEH28
+bZcxe8tbYHHiDDmS1CFlom2kfKJIYGQ60lP9iriAz0hBJTITp+SBJ3zlbt0NDlh0Or6EJm4jMae
S2NRwqlXtHMEO8C/Zvr4cn6tdXZV5vwbkAZZqOzlL2T+SgTPZ1YJC5d05tXzkaRX2zBPLx/xBPPS
fwgB/Qcjak/s9oHBoVjHai3AZJZgIuYSPLGsCRH/QaR/+U5Mxfcf3RALl5cuvDiOobthHk3WUNiE
u8k2vuWGbYCsCWD4c5EA/hW8K2Pu15Nav7AEpjBKU7hRMLDzyM64/r0lrJorMIaj/FAcM8w9zjQE
CQ73282hbMuXPXOTtKeHqyJXzs2T6Vx+DltkGukP8TU7xR0xTJ0stigYPrWrdMfFzRxytCW+lRWA
+1u/OgNSBoGJmpfX4XmlpMYjuSy4Y+9yjs8DDmQPda+GRkqIG6b9bdIRofYN4flcHt4+fKiO+Eeo
GJXuv5UACZiarXQqXg3zqp5K+EgHFKPJ18Tc/LCE6ZDF4GZR8fuxpJsQ+EoU9b5EL8aj37Xk3D9C
a2yPBFUxvOYqA6BLKIhnavkjdfdwDUUnsu1vSksVqzrlrzeZuCnCshnOZjUGAcmdb5P9oRRjo2IF
g1Hiw99kuXTflLW33SrtVenLPSJbnbRgyN8O9M41SkxowNuLWCm2u+7WxTfKjJTGkZzpy64mRQTF
jGA+tjurMHBNZNTwWsPyRbgLpEAXOUNB3R3Da1SaFMF+jkXb5HWFRAg5GHM5gI40c2mXQ/qNTl6N
2wFRhW9Jju7dplR+/CLEag7OH2tprEbD9E4mbnwGPTRX5YHhFN8WUA88GJ3x/TrGK2Rwm4s2TmqD
IOx+gKEfATZXPPjuM7GKy7FyD/IPH5SyNumX8DEHm0YhABOEWnwmdSnowXDCmPSJ6Y8zWiSzyWtK
atjXFmmLnLCBU2wBxW31Wu9bqDbYUfiZSP8aDtGGHLmhnnPgGMPvRIabVNdprpOa1FxMdjxssoai
Bot3aieiDiy6w8rm3HCskWVsnxvIwnJtjJl7GP+MaLqd79V3wzP+QJNCB9XTgN+77RSWFUF+rbtU
MaCHjvzIJ4NiugDKFRJ7vCR95R9OYt6BaoTxGUtvdCc0zWkcrVRWQkybHNWF1LXuB9z1QpCJfcEb
SKQTmx+S6CUKCx6ycQ0Vzru9/R1uElemr91i1CHHpJpk6Y5gaHjJ1OW8mNbgJVphOZvj9nk+iEIb
Y36pIQt0ap600Qr5CzF1mzuQSb5lQnyd4RFZtNsGIQ3U58Ma1BPBVck30nOw0HMG+zwrspIr27lT
2nsy6VH4OFu7Bm0Uvf/zAAvxtsMSzGQuxjklL+4jedOS4GF3LzgrRV9KBUjmI8Ha/eu5DUP19lwT
a/AZSTejsUpglC5mMQaFEqx8/WXSVu7pVazBASAjkhF5WNX5BAlZo5KXF6GIS8ugAX2t+E0CY+eS
zqqbgRj8Whw82pa479I3aNELtNdUtCb5snnAf9WDYc9pX8koSHVeUHq2+FMVUHgDm7xpABu9vxPA
o20yAVTwLRKTnWL9OaH4sxW/to8WWwpymka/i4aPWJRzTy1pnZJDFHy+pUZQIivYmi5Cfh2UGzQd
ecgcauNzJ8AKxtCVCAc7sHhDwmw49oTRglq34C6Qo/YaPMRCHI9kGRO225BdEkJNq+0Jvs6PHcne
xntBMMv9hx/KhgUOhG2i+4qXEGLmTkHilnzkOUrhy29s4r/hMzjTUHdCV6rqcewlDVjGCPK2pAZK
GkluRsdChZG5+yplEfruuwM5FdHvfFzifDv4e87e1Wa30ZBJxbpJQsoXT8KZ/9VYuB7WyDzFwzHx
hQKF8+5giVmZRVJmhpX+HHbRLn4GhmMkLDVum0Iog0KugH1OuK9IEdyDdKpeMJ4gFe9CnM+3YZI4
V1y5QZSuViRf1qTjNxjQXTCa0GNRQhP4uccyR4JlW1ZB1ImiJXgl6DHCq5BxHWFbIlAZxQ4Wm8QO
4ZJhwnnzhRaiCBWnnLut/ExkcxtRo+IQ8y+Nhzq4PMSfLePw5BsgdNDMEOrfC7rD9L4tb5XP1QYN
JVrsMMWOAIS4jfok5fYZD1VIDXem86VmhgAhIjQOPv61ijzXXQKwPEptxUg2sRxnWi7Y5EjHygT1
SPU6u/jO9D6gR91xTi8ECqBnU96Wpxl+PGhgi+XHKiungPsJDqP5C918BxQTnOFDS0V2Pdb+WVWw
mmsFUwzCmfPWXIlx/iEnyCRR4oJvzZ4jN51ArnrQOci6LiUxCZAR1mKlN5/bOy+XGtYrojB/7q8U
XD2latISUr1zVYfYjrkFotCtGODUMyYd0JSSJFNwg5wU8K0Gozo8NelNVl1OL2bufOIAl5U3LbDZ
OTEstw+PmcqLkvvG9Gg4IZfO7pB68UOZpGh9mIy7BbUUCczpdS9b/27EY30oMlPQPtcpSYoca3B8
5t2pIMIiU0frz2U71DSw0XQKyEU2M6hRzdWQ17eV8mLGwWKvQCz4n2huMCdsg7Ee9mfef3OWXZvn
/GdNSNBN+9MZCY2o45Z0ZkfBnp5sr/nHjpOEc3Wy6gCuzr5EJ90EK6oUIp5jjPfjoxr1pSZa/WV5
cQCS7mBFWNjprID8p2nhu3HjppHtjMT1FcTlkoYji8adw8588hwN2cogHH0ftD4vR9GaVxl+xVNZ
kSNV+gR9hxJlUiRT0moqqNxfKZxeEDj7mha+8JY1XwQyaUnxvigwSxeGFanbo54ddValwb/HA350
QZ+cHq/owHVPcaSOdYNReYfFKhwbeEk0iCakETIyB9z1FsXhLvTW1stxlLur6W/OiUwp6LOSabgY
46s4RkHZaWZFtxvGRkiX9UT9r6WbFiAYAmELzj+QTstow1Fmly6hrMSALoUFFy97/a8OdrVPkl7b
lR8yUOqSX/2F9pxHTJGc5Hi+XNhf/wT92ZoPum8IYZbkIlGUxftuEdMVlv52on3+xo4WLnQZMHuo
DHQ082MVWdVr94glf8mEzBk2nsy2Ns8UhEHpBPnmy056ksfUyBEJY0+Vu4ulE4q0oA1Vx6NaSkqq
9EZq2gL/TP319figrkXez2PVkpw11/3sHURlMtkOVILxjoR7LhUkwR36pcl27/02sy9ttkLTKb+o
m61iga3q+PhIifZ02ZPi/2SZ1dWcq7LIsMcDpccWldM8HOgrMoVMzy93jahR+OncdesVmt+3a2MD
59qFCwFNwpap668HdCKk9XDiiAA71vDKZQt3QwDgcSt2xKk3r4OuO/o7eLVNI4dh7p2P/LiAYJBG
d+NapWY35wh3mxqY4U4KO+uD5HBENbfXyocI8cjDIsTekmHmvm3h63iEDGAnxfa71DS4/mTUiFLU
ma61bQVPyRTG1PmPh6F5qIgJctaA45oB48laUPO57blFl6NqsJaDm46CIvL68X5X2fArGgPDKlM1
C3Sh7qZ0IgrteCwKOrUNqtd30Xtq1SHZnv3RVe1PPyQ51OyPQiGJD7omfDipxqtSf2iZdRu2uzOM
VzyREisCOro1FD1QcqFmFoxuAiXh4LFQcFTVj8GhkMydm34xZuwnwTjrWAPWKbCCnb51itwoLGXs
kM8Lgz7dPhQlyHNUN/ZSiij0WFuUn2tJi21hoX2ODl207wPq/82+pDVbvjiWTFKNnYbGslpajMIE
8syyJEdlMwfxjlnhNyZ0NDoM13hzmS80c0XxR9D7i2s0VJNP7hyfu+A0jLOS1b0ohVGh70U5sN4c
PgJpaXJq3dUGBHa3pU7du7j+J+5PAchzuFO719uB0CGv/2EA6DuBhmFuotAohd1LUGwZmmkPdAHH
ssKq7RYTYGr5E0cTLZCb8uRsHjqK0xuxhJ6THQLh5G7WsoTcoo/1wjWWprQ9lpNLc+TVI8u5jRN7
h9osGY7DujRAijzPmqo5VW4snTBpdmBPpkEjiK3m7iW8JUh+LlHX5t14Pk5sExcCuZD/s0kMXo7f
fpzdKOqOxwNm9BrlRBjdB7Cc+LQ1TUQsY+vcpFkOG15PNG4UwlDP207MdtCxGCm46Thj7M/Z0JaU
J3wGnkhp3iUPtaURX343G6+TcN5DvycQEpqbjwIsYpXhMwR+lgshznMKRpMl7IRJKcTgRuOY0h70
QEj0pWylhSjJBk5lq/Plx5BCWN+4cXpJ2cnM4caHZIA575jCEr/fplmj5DObjrrJiaTBkR578FM6
+CeI3laoDhXlbRA/qa7eiC/2+qpfzRfjq1HqrRbdfo4i/hMrx/V95VCXRmkwZJm6bcdUHGM4PdgY
588Q91eZr6GMDWUADCffEJfS/aSxMWb1UD39jcgCFup10SIBmNJX+5wT1Gi4GvCBE1fBxvhX7D/a
6lPK97giwQEMCL1aUMDOGeMhXROaWK1em+XCpet2BlJfEB1y5qzMgWKW5LIXREuqmmPLGr6W1fat
uQpR6NjyaFVsL/eqrUwZcxoe4SY5lj83cFEqJ9a1ynpNd7mGeIv1C0MCDBRrmKlVHBExEnz8hoqS
5pvZpkLlimVd4lMBWJl7irMSH8ySohbK7Gu3eX+BDvMOA9qLuUCEI1esrYrwF2pror7MsJlibwaF
L/zXlgO4u2C41JmrlwJxStv3NnwsYHO/AlVnDyHXDBjA/gNgmoEZCz3jgho6UAACkRybjSZOrYZ/
PyrSaocNVCKh40SUpC4IcRdwixiGqOZoPl4U8lNCAcavfypV7tOiqzC3EHK+pSKDW/ynIYgVy5Tx
DhNMLp0O7kUxDaFsnoUjLsFbdDGWYcGmbfAs7qGvL52LXrhQvEZWHnQvxmRpJzeJeLB226m19vaC
HgP0Bt0GRh9uobdbc/HPlrcR8csZzxAI4OQDDXn6vGK8r/+zus+KqSJxz2jE74J5BNilaq6OvrJ+
EGCPXjtcUJpOpU45AVQ1BgwFF3/XUem5Mf3f3eqWeJEd0F+B5Z8ga7nejZNXdjBtNQCTtxaV4uBv
rfYJrfauXeOlBL1jYhzxqrvQ5BaST88xJxJlgkKCT64DUioP1k0jwcxD/04jbMQN/Y973IQKVs4g
hIBlrcPt16D+jV/JfJ9wKJQHvvh+EF20c5YwUWYqeDJSt29JmD+IQeed+4kVIpB7pCV/yZALNkdS
Ogg4M2YUkmtrXMrWMcwek5c1ju6Ewidv9w39oT/jhA/4Jb27HvF+AAxCfQESIDoak+DKLhRRSnDt
yWEnzliUE8iLVahbsYdjTK4VF3ZtrzMRrphRqOnYwpT+RUVUBv2dC69Kc37872va6yR6LUf1ZBk6
9HBPTQuPwiRceLZM8PISvK2Pj2PLsXHQicHP0kIFyDdwlSQnyqa1Z9uoTFhP0qawVBQP4y6co2Nc
TfenyU993PAYKghVTXCaODbFaVHGjpBBSMz4LRUtvK3MQqKaJvUuKzAmEuSitGV1649p9qokj71S
7SM26GYC2uiwEpoVXkGLsfOfgND6+S5clmAxXDhxBgaULxTi28LLROJIRdkBG++J7mHP2rY5amHf
nJwfilRF3pTIOv398CAkDYZB5UU/PzDIh1Y96/FFdWzbof+FonDCiNf7vqB5zMXdwGj02BWcywGO
o5pyn3wAEjRi5Jhav/+OnEZYLa0o+gRITX+G7ckw8548DbxOPK1kNpIOIQBFwcEDJgzKElVjjfK1
6w+DpfjaqJA2GwJVYP+u6rgyWyQvpwqGn7yW/haKK7XDH1JbSkYZovxWwZ0nlVIqchg+bw8iqLQ+
z0q1rs6DtbyDrE7IwumNBYqaFEmK/PnR2pPxY0nDZBdHPuR895edo+e0saPAoqOASuZmvO0vHmh3
oyKtrL/VzQ+RuDkGnQLEczVKHHbRd5pjNkCu/NOx8pwVWstm1beInxcH0RY5woB/GM8pLiSkhVij
8JTW4dPEruDZPqtePgA7unwqnD/L4FJwyO0YNR5c7KejT/WkxUfMGOJL1xv/NClvzo27/2XgNbFF
4n0mr1whNRuXwfoEvqT/e8QSxJx5tp4uEAMe9AhW29U58qhffzWUXt2c1mCskBRTri3E8r4hb8ng
57GsJlyNEXMcVW5P2rV+vg5ZxIHDC9dfQEP9Mz173R24EjzhpDKzEi0kj6ES7JGdsb5s13vdPVr/
P7otqGyTw6WocGgf3jOr5yYpj8vIFv9IVtvSZ/TWagl9nBh0yyv6djaX6FpxxKfAOhEqMZ0EiJdc
mXil6uOVVYT43rtKEgybUVdUBP3lROi1iDY7lGO0JFKvoUxEf/2S3yoR70TfrqI5Zv7z0brIQp6t
G6LvYvuH+yfG4m8lqddIRN9a3jBGzYt5duLrRjNBiAV4W8Dr0M7nZfS004o6ltpLodXXor1NA6BQ
8mWf6HI36Jc9EYVfbnIKGOatSyV3zl/GgFCe+9qO8YnDODEvPnbp8fKX9tSyaINf7GivWirHPn93
KwLesFMICW13zG6LlvUkQTGvwFTUND91Ydkfv7qwFNCCBmHCuhF+GBF7AqDhI9Z/efx+ggMdAWs1
rESTcqndYje8AtLx7xf3NdJVHRatEFKPPoN5tgMI2kGYT3CrTEBc5bz3N8WvStduISzn9/3A9Mu5
/8iiy4ulW8ZCN18Cf4JOq3/UrJEhHKxiGrzpxsZzggY94s2ETTEfIGPhSNefka7iTYrT+oASdlkz
vW1UxfOamjfMIGLTxQ9N1vMEi2DU4798iQNCoM+enP7ki0Eyg6jXiCQU6Rcne/U5Q0IiwPdaNOLf
7+aAWN96FfGMhbsmCXeTl3tV7G9o5XXtnPKqlwhhuwM28fFT574ggxGz427TmUy4dp03RHsIr6Wa
h1YsmE1oMpSuUBd+WWeFoj6IuGuxsbBp6fGu2L1DhJ8qD3vZ1rHUpS7/36s7QkdMl9CJtiHIhEUj
aVxAb8AmXhjX9ic/CTCXv5VrzRVZ515ZmdfL72Wq9Wo1b3kSHjlHTSQLqWgOeNiBOWcH8hYWUxZi
zhnJXi2g0TyzLsex+d0hcfB8Fx53L/jpiIPsnB9mAjdLanJq8RHIVmqnHvPLZqsxU+GvPoVezc28
9GA08iuM1zGqTjO0elJPuQf77HaOrnzFieU11iONiMErmzCZBKW+Hvfhx0ybCsLq4jKlKfNnqCVX
Y0cW9phB4KPNybV+ABd38V0FDFkpIciF/ma53T5ypF2dzOlUVufhRCBWZ6Z5pytm7moT+hxK2+19
t8PaRJqrLbbAd97NtBUsEGHjqLPkoHEkQMaqG3szCiZ01dloWuldahoUSr4RnZJe+VWUP+ZzmFqx
ExStI8CJb0aji3ZV0PwV2MXiDLq0Bh+qrXMYSciHg1I73KbxdvTYskAN2Eboois2aysqmXACGLmv
zQm+K2DUMUvresy6fkwk+CyIyOBwvopr1tkrZcubWuC70dvHY64tg/CGgb1FXfjltIN3iLNqli+Y
EKTG23FxKnBi1DNE6uiXeBccOYQNx5apvg5lhXCEhKmoCX1OdoM2oA5V0epNrijXAlGFhDMd3e5J
NbUov8QjTZQZZiVYi0z1FbJCLLOi9XxFdqO18NPuEBw2Pf1V/uosp1nYFUd7lVVl2oHZccyRtHuC
0ktVv0sLFKQX1JPNS0+Gu4101cETUvt2fW4B7QIkbbtXA1fJX/AIxMnlx2JT9Aujn/2x+GLBDVRU
MGB6QmfZZ+VDNasTAluRKdoa4zkGLJn8RC4SlOG5gH53utgDUegjHclIkVGYXO9DW2njW4UNtr0J
msGQ/VD2dKJCu/NCNbrnopxBhsi2F+8D5U+4i3ngltlY0lxdYWs5cfiOqYHpUoKtTpIYWivIrtRK
xsNm47UtaAJTT7bknQVantXV2FSBo+eVpydKbcluDonI2gYeQtioIYDASJ7i5MK+Sqs8A/Hg6ybh
EaGhg4RiAyOb/ZsLH8j94XM4Y+Is1A8ZlKSynvxLCbJmiAcV/T/5dBh00rdJLQBzzfF5DefOSHeL
zlry6qFNqtDRAIOiWCfWV1Ehd5gSbRVIW5LYtJY1j5g+oPHwx+a8/MDeTyDXwENyVwoV0dy/xcVK
4oEDYszpNT3BogYPOD9O5QQDMVRnfa0cnWezvzbjGxuKkxBDETb4O8nIiCJ1Hjzxwg+SXTnJcxLm
FCYb0qp/x2fjSwGidHPdWhPBj2PHpKGkoymCIJbTiGTS+oBxrCErI5dMmvTcUKXE3MDivRQSLtWq
V3+RDOY09tHFbDPk5bOC4FKspA0BXbEw0HsV4FG5rI5RXLPhAImx6Ul0OHUW28RKPw9duZocDR8n
OycoyR7OsS12agkjv/DsY/k83I8rOom4IHOOpVA1yVUA/gqyARIDRt51lRUbNF+AiLROUWytQ9c7
yPFXMyHwnz4Jth0JE3+/AbKHihIZJubYuQWDUmRr71p+MExfOO+PlUomjWaPE/jQpOiEV8ezjyFI
23JvWgqDF+EQzBch5rjbk92qfyKxBVzP+PRDpOA2CJyq4DZbj4Fr4xMOOaDnmYokP3KSMJyWD6Xd
87dWePkDfe8kaAoYqyTySJBje9g3B29sdGiwNsv+P0tpQNxJS+pk7nbP8Jpi2UFuG1dqJeLIlfPH
mHEkbsr9Vsh0ZaSDNRCS11v+8AleiOi74FDzPDycYNQkChEsJcrYfwtbn6KmUGw88JfQfGThjEiM
Tb8Xx1bhz3+ZMIjnCQqyPXOsLR7VX3rH0hnXp+THFwIuUNlq+1397gVH+LGu427D+my6Q4k/XCVs
e2icfn9QeFaK6xd//o+2pB7hkQf5JXUpfRQgwrknvCztOHrVV/6Gh6QdZRL4q0dVSjw1P5OR64y7
CFeJRHvBETD6eIOuTkiCQSJJoGhxghIZ0scrio4nxiLl332gO3MrIucLQDo1Nn4cH4xgRULV2TZ9
K2bqvHgrwp4UJenpECnDFeURF0no1Gc9udMm7KhlQImARKniLYhGIdMIOjTRwZ/kal22xXs4PRyu
w2ekJ5yBag3NHFSafkxTkdxmBx93hhRaWZqD7jBgMEdTMdzEo7UyS9t1Wql08ngFa7lnMnhvucWI
IgQCgvdD94OLW4jqSEavpB+PrI6JDnuf5D2QozH34p74jefwtLXJvqsQKWpYDjbbnaOAjcT/Sd6y
oEnOpiT7w5czhumKWA9UCDQX1Fub6uJfJZJMVCh0Wpb0p/u3tHvZpvfQ7bC3gQFwBf1v7wUlS7rx
ccZKdv2QaAeOUndjt1ghD+kqGEnLtyNjwZOsoCebSWhW9LwxgXtAnMre3SJxLpyHZV29khk+U6YB
VTsRpwOhdzUzZHJhr+ykWvSbFRDHUHuX0rvdp5O1jsqLvbD6IE+DDKiG6RN5xxBcoAT34nUlxYnA
r4dm1w34cyQcfsNTbRYERLnelllEOiOHGe/kWW3FGaTJOwonmUsuo5lFlXk1TlywIQdq9mxmay17
ruMRT1315ZJyhNU3cKzoEIfC4Fm2VVuL0EZhpcaFqcjprfuUa2/LmFK0fPlzMsPIghgMwVx6PD/9
sZ52cLGEwu5PbqSymUwo3B4yNCjNZ6Vv1eFw8GCYp2Zhe/kx/hRLWJUhYynu0d6Xt+3LqgKTnWRg
X+lxl1P99xjXdjQB5Ktfrdyj29LxdjF/IhexYfZVjb8tzyqpAlUpJJi0GGVRh6kMQ9cydm98sIVh
UlEKVKi/RkXvD1JMh8NDUv9uWPheApw1qtbhVFVGNV8seobw4TvX/3dsl8ptHfwIEvlOcsSifVEf
Taz899dC3dxCRK+9vF9KLE5Rvt7Fu6UMjjQRH9rSkW+z38dpz9RFo/RoiJqrFn+tH4e/xocY96b+
uF/7FC2MQSJJ5DX+GKdZToeCw1Rsvd7OA4saK9sOTEZvAv/TJgwLDMOkrdeMLn7WEjkPyEnkH/fO
ymKTQfX7+q2LbF/9UK5mT7c6vA2r0AJ4B6anRyd5YWWu6RiG44vJ+UOdhKOufknuRQLxZ+WbHTq7
lUHAe9emFU8+ya0GopQhFfbLgmOSIiteAcx0X2oTvBBqnKhEnL5Ke9Hi9oTUqImJ4LGZNYhfFZJY
l6NqooN4yptAnq1+0lgEnJMmvpHvw3b+J60gpNb2Ei5tpN+kDQ6egntR663YXhcm3O3pqA+NlrEd
q6Y+qzXKxUMxZEEKwDbiAmLqORWCAFqLZwhawCiNPeg+BVPmHHP5QCnNiqgWZLWGeMDpld3hsDRP
uvJVwKMbIi3E+iQxLKXwMACh26L6qRMyuFJEno13bP0tpvYv6QGFhV3pSyOiLNgO9wkd+Xmf4msQ
RNRBpyr3g6rQLMasFMm139mZYUTmg6WCd2rQZDCobLBi0cMf3JOhnSHV7EwD30EMEg7NcbX7s9IM
Bn3ZHxwunZyt2bJZ4nZ+s0Wd/7IcdzzS23H18wuizf7HEn2c6Hlo9NwFvTuSYAL3M36AWldf3487
aBWvYd6JgtWfJXy98jOza4xIrIjeE5OOPzJtOgFyN4BY9fImCjuLesi9DIu97W5JDduCUbGy55o4
YyiykcxOBj2kfceb9vw9JygNJrqRZx0sEwy8YEaN48jf1qZhSE8Ie938tYKij37jrzuyed9RIf1X
7BiP4wyIysyzZEsUg0IkO+cmnJiUJncQFWOfG4fQ9KrkzY7YIGDNJFJAtMwDMCPn2PKem36GGj2Q
lTh9kuXWEuo4L2oWcDXKH92vvqiM3Dh5EEevHrXx6Huy6JnqBU4iC4cOzNrQH6HmxENv8fBfoZOc
0lvJ2MhDKAkS5p97QoxSiXRvyog03ItgYg9Uu5g/UyDbvS3ATdIVhV0wM/qY8Q2R7Nkra4/ub+L7
j2Jyk3LcERdiBcbQtSAs+/hdH/KSvqbqe2XvulaDAitCOfg6ajab/hLTxi6kJ3nmDhcKdeDs7cVG
w3aGPAlFEhsXysyLE84HzUFqZGJyT8SYthQmqhNf9d8Dq/tayCuw6fsQkDfLkVFDlxtC9u+4VDqZ
efxwWOhbt+7UmK5lnHZBa2mSN6kHjRiNgNwf847ylqEFjpUfVn7w8HBWOo43gIou/2RNg/2bfrhQ
SXBrL0u/giehZuFF1DefMnb8zlfXfMqT4r29JKbgWKwWv8vjOtEGc0sabLOLSJ7XB+t+ZS6igYWb
pWXNUjzPHnwFoSz3BsHkvIb3XxCav1PVy/GMB7p+wQBPpzdwDl29JfBK9CRUg5IvUM7M2LQHkWyk
P0T0676EMI5xG5SJ870NaLu7gVWfq0xBxdUey83czJeF5y2W+8xHJGHilT621oRgj7dSKdAf+ZV/
vjbsEyxyvmJ7kQF3raXwpRUM/xbZcQv1Nj8HzgxoQKoGssVS68UVYd/++5kkM5H42gMf1ogE97qR
xnZvHPvDSnNKOlZ5cbf7hzaiQ1h5vjAPyqSYJMW3mEeUy1FhnpagtATmjwDp0g/wjVpgMHu5r7uc
d1BpAfBCsqNF3xUP9OW7kEd5X6nqJoYe8ou6JwZCcXoySqHjOdw8B97upTFb+uBtLTJe7SlfgYYO
emZ1qcxXgdDYoQRsceeOVHfsx96LsrRNcMXJ0zBvQ8LbQhTR2rnAzq7824trk3e70Up4LAz6GEn1
acC4KTyZsaN1D6lzUkfn0x04c6VKlGoGOOD9i7B5QIT7FtseHn3O9tZh1fi5yz8rYI+qZ+wL0k4a
xgbR9GJwi8WYa4H/YM+dEzRU4CRKCwv5BFUK5v6h7AcOlnTQiLz/hABk7RyfIJ8Ia5s0tXpCdm7k
6vqE9WDbPHrI3YZrzAw4JxcXcbSRGzV8QHU6fiPtiqTHpj2QXytFimbGU7DtgMt3DsRQBxXx4FNM
lrLhPzvQhnYD4sOmVV5I210wDLDpTHCmM/Cax8qc7h4oMnTt6N/b9o4An8jvmdyWvLni4l9JClN9
Zp8WAt3/djNWqxGAkX8bHwa5x9tQH8M5E55nrg+UZlpjg/f6UBvAbw7/p/n1BXu1WUS7/y9OPGqJ
P3XudNbRmrPu8GGQB7SATfqa/1yue/kyN9env57tNtzEJ+CRlTxzyAk6EIa5mN9K/99nFqeiSNoI
M5HMTAI2zqFH3g7/zHHDTmKtI/Yzan+w+lgQNHHs7DALP4/niaEBzE4gphdPG9Pq/WG0crvWXJDg
JY4t9Q79vL0Z08ko3QSYOlxHFXNpLIJcz6yOuDmqmVV9dAL9dJrIJo4icmFangZCz6pOOBNuLUxP
xFYWzcao3zBXLprbGlgfx1r++cSI/p+UhjjIJMCoGlL1cFqgHI2BZMsgOssm7uue+3YEtBPds6tc
rYN4xAhRF35CMN+uh8fRibsmshn/qiepc5aPuFoRJ51VXomJfHAQsuaa9KBOb1IB6CD2JJui/Qur
DupFJTnh0a+rfHDhQGFDbfTq/EEj7pZ1mTw59/LlTiHqymWWtCuvAfNguUBqhuZU2kOuKHSlB/CX
xdOqi9dX2OwS1+d+7ZVoPxFj1rEdddmfNUkKqOHra/Vhl7OWLGtUlTkomAj4nvNDEUcVtpyeBU5S
L7//uVY2b0tvbiUReGqFktCxg3uXkRpazSLna4t/9SWFeq6CISlSsI4KCQRxoZq2ormEGsJnH80d
9rAWe63o62yk9LOgUg6n/sYQgpHmEGro9o1wq0cYIbhskpLQ+/s1R1eUh/cpU3lMaPpE52fP/qtO
9wDy3j5Fa+CH90/PC93XlakU/8/9S/KCRxNMx98H8FCALwyucIQh7gh8knYoEg/5t8tE4aOUwRxA
T5+V4g3NUGwJf/vygp/sH/+31LbiJM9bk2gc4G2OwcAcdbcaEnyD6kXQpx9CxUzUrMfyjZfxQG8d
jjecErb82v/Dtnyd81I4wMEE86rmbieGL1hGwafVF4byrV3XCyRZxf+YL1Du4Z4geyZeSXY9Ah2x
v8VM5rsd+btKh5knclqimIlW1SXxzmjXXOiijG0Uzzg62ntd6bOYq/WY6v7oZ3VcjBDr8cF0U+Yt
HzAjpCG51eH9W+0l4CYsgQOAP3969cDkK3E9AteV1n3eAzh7h2GVk0svaNcItFsPpQ++HKtoJMYo
qf93+WGKEtLVX9puv4km9oXcmhRLohvsg4Yp6S0PkYEx6MSOOzHHUEceJafa2tuWew6Fruyrh2mL
1Gz6EaOeZ9ENB9+MPg1DdoMi3QMoOJn6sWwT95NcUXhvt15MCsEpaxl6N8gsFOqE74gmjtUpeMut
1DsFdTLlWUPZa5SuPE/g+96u/xwpUNqu+MMBtZ5axtmX5hmpEXWy8jEeNT+5gDoZMNJVZzna+Pz/
jUja6qP/eERsLCgW8gKmIQXY6eLBsL6dsBNhtEEjPXQMycjpXoeyDtx3zaTLF7zvDviUSV09p1VI
FXrfQ+Bsde/jzcAGILNg0SuoH1Tho/qaeI0TWHpwcL3uLSurhNocW6LI4Eu7Owm1aQYL2tZ7Gn5B
5iFYCSS2mUumVx8ts8ESuMWAUlWq8jLnRNp/bQNlO5Ja4PRvsOJo2MVl7KG87tVnGSCtSU23ycft
gc3TkmEWkl5XP7jDljLHSXfCgfSbgXhLNFpa7L0zPEAY63xBOCUrhwvNe7uCfwQaoz2omy3kPo1u
lEcHiXR38zJRJKE4aV+a94tp28KagIeoiPYC6Mt4VheS4hVjLoczuXxC43k4uXouu1/NQKjn8RdD
5eIVLUes7NkPfob7TZMwafm44L1OV2OlO6aMosiJcQmazrY4rOTTJ+5menYDFjroyDzREEw9+gMq
vE+TXOTv2sHiqNoQTOIdNHvF/0iN8OhPlV0X1hAOiEy0Q4hp8DNjL5HqgpX0RFk+1mhQuVCEFUg8
aCwLqzGCaZ64vKuUwetTjqwTjS43ci9xHk8r/lX5C3bK2wNMh+tFKt2y9YtZ4je9F+RWUFqOVk75
dJ+PMOijS3Rbzto3Gc2OoavRFyxIubgTgIsp/ZMbrCLfxO0ZhqElGyZBW9GNbczQTRaqARwy4kb4
LFPUqLE6PZmrExpnpsaFKg26BZ9TV9OVZ7+pAfCngbqVHC3Zp4vXkLd2Jd0OISjNcQAWDv4qDGn5
Y/s4z6jzpBqqm/KFKOU6kc74BSG53Wqs5c3DQvdymZvVY+DttRE40+p3+VG5tTurp/0NeAJG//yD
+OiFCNx3JfkF42P3UA7SCxIEoRO9NrjLks7Q+n2+0rcxpRwH41HRcPL1f54RG1lQePlBAWS0P9tp
Ek86DNWMq20xN2WioE40cl6Kr/+B1Qx/hMfFw6vx8Sa66XrqrHpmMDujfW8xIFgUlmLkzvw0LC/1
KITIzqDDHFIBUp2pEbkNXaAfF5+rZN9xE72Z5LgB/xi+WEiUD1QvBRCQhljouhaermbgpbf4FSdi
JjIDKXe+ZvBHuixJCfwfDa2JpA4ZmNvHP3FjaypM/kt3XzGgKstWJS8A1xzgpPGDfQZQCiO9D0M0
ps23gvMijO4E+86/W5W2kANLq5k0DGbTYZ89489sIl3O5VKjXbFL4/Q5RLWqmRHfs/F2slBh1IP9
EsWv/pjWrej0E4x/sP7XUvbrUtiFPcQO5oFHYdIdnu5ps2ZP9OjmysWy2yIjtJJsNs4jxGhMQjtB
IOKqgKEyKoN+JTVy4KZOEcnLJoXdWNs8qKvouHB4RQzjyqLcSJPUwvzFlai6aIc5om+LkrUlowyP
FCNUTJWkjPU9Z4o88QcvgE9H5mw5Kj5maqHUcrXDTcOMtukycr/7d8rH3+i1Og9uAzXB38Pbo5//
AVja1xNNPgN5ejTd9QYr0UwGOPUR1ZeXnh0UEA5r5evFdwR2J5YbvjU2QaitjgzE3yxC3qOjDj/z
y9Zs6x6Xas/AZOpFdra42G9XjeZ/EpkNSqo52ct8YZ8j95mFQ3fDkrxrsluWKApvZ+dEKqv9YVJA
rUcFQyo0Onb1yLnQBADMTY10XqLznSeue7+Udkka3YmF+yDUwN/dSouj3li3OOMZqh+8sYOacv1o
E/DRKBkiWtp2xr6q4WnS5BVh5+aBl6z4br7SBY9aS94l7iPZ9Cws2PZkIH5SVzEH3vTjvSgu1LW9
3uoc8h/2Y8KkD4b8+exWP4qSwq4pr5H5PIEqp8ibehOxJmSapyPcyYbB7XRA86J6lqEKpBezMusu
dXiTVNQsk/USrERMp7ofCQ69pcHVhwlBEVhfrC2/SnH/41gZZG2kSaLq6tCXquGmoEPBmsMIzThD
ZHBnjsVDyvUhFtRsRHw2c3OKib5FP9OdOW4hdL0aSuO/foVxyRoi5osttDVS6CU1y9PIJ4TOCWW8
PXpec2z90oU7zpyUeszs3zpAZWXgV6pFowjcCshk/30zSv5leb2T7otlTG2KyHywLJHhKjrHqWwE
PeuOmQDzpjXqcfBA+H3cQqufb6fC7k3sXP3GoAkN4S8qu+OUHT2kkXYvl+KBksGBoxNKd2DDDC2w
aiJGCp12AAv+ZYBsKNtm6+HI9pIor4R54h50sgWJjJ4/HcMFecNpQPaMEswO2U4HOsbUVqnML07h
DzupZVAlmGMw1kwRCZjbeqL2eeH+F3ag1SarUg3beGGeiOwM1E96kbtSxzkZUc5dqwPQLZ9qUtp/
8xn3sSeH/RGgycwY2OU1FiQj6lVhosZSrPwjOEP4HaAddqXkzjc85nUDFJ3AmeAUFqNURiVk2wwu
HhxP3yAmNmVe9cGSGECjsP9aJG+SdCeWLghOaTPXqMCYfUHYpT/7+qMX3rMlUWSYqmqF/Sp6MrVo
pPhRh2HCeSyr45OWqWh5jla37bRzROwgaSL2U6pxCJ8zzWRAgTXk4Bdrn5lbwBGMvpDabq6bc8XM
GtsRq7ermYdepr2tFTxIwQD+q+7M8eAYm4Ig6DP8E9bsLnNFO40q7+ABdwC/dbpL5K5St5P4vhao
heu3IuB5ACsW4Ot2HpKfetsoM1zm3EsMad+QHQGDv0+KU2FKry1nZQ1/9daxNizepNa7BtOh6S19
CqEBnfehxpPsNNBijoYJ/2cbjtd8UX13uedOSQTp3NCzL4JfVlPUjGQVLgzABLf2cCe5M/Ihx5aj
kBgcss5RGbQqB5lkWuOPfwvW4ujY8BYyIauNDukPLfEI61HuzVIPEQpcVfn5NDoH/S8EEZP5P6Yi
fNuqA77BBGcZ7HmLws41m+W98FAU4TZK3jEqmbotYpJUluBTpZNGm5HKzJA2BuLmPG3r78cNJ2HY
w4O9jUvATpRRX4M3RFAdL8qODLXXxSF0K6q+scubs97mLT/FdMjL3VhjeWFsFlk1cKaGSEFgG604
L+ITwmqf9KKdfIGdBz/i4siVSqpOFNkwBYR25imuKIO7/cHvxuaHBXP/BKU6lDtpQfUJHHi9d/Dc
E++ZO1u7RPkSgFf5/DoQ/gm8dPlYrhE8CttQ2qlgBFXAmVHoytK5diT92fgFNy5Xkgw14jOMOJxu
WsmdV7BvsETyjf42qxhRHIvoirj/lZQjYAOR9kWUiD+cEmIBncFhIrBzr88n5pb1T4lwbBN4FJdm
8rDFR0sXGfVUIZw2xf99qk1M7p3vTiwkfVHJyOY1gX1dSYJcbb5FQ2O18KtQLnJHeCRPcvX23DHh
KeEm2TMtGSkQnZZPjq5/IGMyIAZWUNeps1gp/4JO251sB2uijYQEwn8gkqyAlF3zNTzNykMDXJ1a
6E7XrVCCYvuiShCgjXNlU6EAw/jKBJgJFdmX09IuHYM5xlD+OHNd2aVvwADdLDB66FYZ3qKpQi95
v4KqJqygiAexdrK1fS0GqXANd2ltCDbkkUEYSOlMfX6wa7E50yqzjC2JuGWHRsK/XI7AyI4EvC4h
zp515Yykgjfy3WcDmA0hr+TR5RGh9Y4/BvA7/Wts7H9VILBw0X+4Xus+m4aYvhc3PXe9uE7HHli6
KoDkKsQHCyBHTuIKjTWMxHyyBV++NpCUeANSu57ga9M9R9AxgdViRGNyOVxv6iDdODwwY13RSViT
9dBfg4eeE5AxtrACXjEOjrwAbd1hO/YxIsYGtUgzs1MurQsrz9WinfhFPy1vgFfIZitLPe9jsmG+
9eC91ubPK9R3IlNxVvPJau7hDMTZwoFhhPIerSPKT3xAo67YJ3Gc4/30KZQ/5fgHDvMBTv4eY77a
9PG+q4lkWYY6rs+wOpjfqEChlPdkpY9EIibBrjSdfXHASahqIFdGrpOHpBQ1nZTD9mZrg3o6ewLM
I2jurDYCgNutjkciupgDstOwz1OSRWWKu4yaJw9zzCSZtgKABV7e7sNcbKlxuo3W5Mcf9qEELEbf
kmW5gL7+K5h/B50OKdjPn65+zc0xUCWcgCU3DiThjHA07oKO269Xq3m9QsS3avqrfLW+B8eq0Hvf
B9HrExPYzedie+2xx093hMit12F2gdgoq05Kkr//MxUZGVSfpUMlRdOGpnN8VnRPmTvcbi5IGGVC
iUm4iUucSTz2BPzLdDe/Is65O5ukzG24Har/FWYXKv5+5leeVfm9KADY7dorD9ACtt1PndjjJhF9
S784WMVWfhFnuYnfvAJziw4OHL8bneamEVhLSL4EBpzp5SSpj9LCgkFpTmtjas3wvyrlT5ho6FDk
3cZC0H+EXITHeeLCDgj9EH7xbwyPYYGo6kr6UykLlHyMVNOcboNf/C0WS/311h8BpC3iGsYYZg8A
6buKHVbd5kAUhaxMFCUqphQ0UscBEvNAzy/JShWH3Sh5rMFIlDPr99t8dh6fgP5I088QlZLY4UVr
EX3TGCRZsiVVJi/NPBYf6mnjle9UxJsa/zD8KNtY2h+jbI/9S7pEEm3uY29wmAOcSiKe51YnfG4q
kAdyOGoqIzm3fE2VOOztlDJOKABNCVa/OknP9uLQZEa+UO2oi/v7xXdMXA8ahHz5o3jMRYPfD9Nx
gqXOxnQqLUXLPdvSEecxjHGZxvi/Tg/EF1fjDiZNzJXPEpoN+Wd4Yh2u+b6ajW76E5oN2zkgb1OZ
ufID7QMFICSk7YR4RKdqkMXvwTWcLOxiDqYBFBIWr+saxhJW3sx/A/RSMgvDwmhX7cXpWucK0EF5
zOqxNPDkoOHBykrVZh78SkiAwuaCHcK6wNvgb7/onDcO2PyXqnFsVqhc+8ykiJM6ujZVsP6MWPy2
q3onNqyL28pcgADPjy/dS7Z2VFU1F9T4KfB3/Eqj6AzdzEnpOa/RVnbJFvkErr6N6CVMUTDOzOpN
KBMzujTEwFRB6eZBFMNRiqTtFMnMbbZ71c/6i6qz7koUyt1uMWmFjIhkFjYV2xc1S5vtdot2bgSN
ZnJqxR9S/H8qL9giAWx114eLw4ezoE8XwCh0mGcx0dVJfro/Y77lG8lja7MArdTDdhJtFsTytO1+
SGd1uVKUonBwriTBFgi5M5hq26qUz9qu/RArN1U8SEUI8LxbZ8T6q3VAqhfhX9z5mRUy4jgnV9ri
XI8VMic4BsJWTO+7aI1FjCNXZ2jW27y+y+4ZT8yruNm1m37IdqrCv+wevruMwGR4OML/Hg8s5w2o
sTsFNZiV4c+Y5dpV4VCow4WhZtUXZI1CGZSPZ0KNC9XtBrpP4V7qA+RNgX+ecKJZ2pCo5Dqr7QIa
q9u4U4m4jn37V3hDjJ9RJ/uOXf1p5Gey+ctqum0EKu3RtlMjkUEJ5T+3YYWHvFn8y3X765riwM6p
tCp68DhND76gqLmhgibcjFTU3loxxe00VrdN1J1d7SN+4W/tBhJfDn1hLFmGKscY7rKz4bapvmzs
EOHnhHuozNkYTQ2YlKoUZJvAIYI3VFtFKdWJv5wU3Ph70XjAGAopTt+vz8oqE5KH6iEYejhhsE9c
k83NHCLEs4P/Gkq8LJUwwLfjntGwAryABkkS5psg/H3vTTt4h5hPxjxreMeIBJ2ILvXWMEevhAi6
WWi0sl8Hx/1qj1eBvl0nD56qMRn0aViOX9FlTGAUbZK8Rws9G7WNbCiog3utsuoUa2JQTFg4dDxa
hAADdY42t17BIOsZif1TW0/g8x+BSS+0eR/afqcUWPnAsQgkYdDaeH/NuvUgpZVAMSI0G7QzLClT
m5G1p2YM8PQo7mccqhCAHDdQGJUKWxZjYN5+dUO7CL/mzwcVPZNz/f+f7pgpwOHTVSdOn27XakQG
uamlyW9KsMqikS4aYG3/mKAX7deHrpnwwDL1uVhdA9HfFUtFzYb62OPrJpw2ZAJ0MBf66HClYmvk
kSp/VKpxgaZhGf/7AyBBrBSUtiQdl46YcrOvG66jqvutjCk9z8H/X165BWVJVOAZof6quxjnWjlW
wMS/8oWQ4AnWgpsoktCJ2g+shq5xGPt8GSNnAVZKWg+pXJPMHIhD4OuacL/Fxz1v5YCz1EDsQ/qY
yJxqMgGwjSsBjJO1ttbXrifxrKpZ5BcHPBoHPMZjFXwKrimsLkKSiO7ZT+2NNURHDjxWCCHw+mgq
p7jpAkgDa3QRt0ftIaPCdeywTaNXDUT6fvGqxtSnj6VtlXaaE6DKTUqt+BULihM8NxNGnfcnDnCb
QznXwDR7ssKVeBG33b3IIA8bBydn/ZutzQfbNdinbHk8vyCiT9nV4YUJzXdPvCSlgCi3Jbnbl7rA
DlSdDFf4IxnNgiGusVCagPCgJyh0hXl8M1JndNOPpY+X3PEORbAWD3toMA5Timbo95KM0T2jgj/B
m1vqK7DcdCDJSyLRNzQ/IEQTT9u2KbGWn/0zz9/3yfgC8v/gLrnLRSNQhvwnXGCxEAkD8g27b8es
zO6B9nCZz9YrfyRR99MkSEQwcARpqiy/xBUR24rFkqvCAK9cVrf+at5gvRBISD8dHNJwuQ5bDkEv
jwZ1gDImu+/qiR22MFNj92ENXVjHEz8t7z/YdUzWgo+UFUovP5L5Ei6s8eP4vOyNIafYI5zHBMU9
iY13Hxjn1vVmgBN0kOwBfJFo/GSp2bIf48mBFBqXPALlBWBla9Zsr/fGIkc09CYMt7VJOswfcx+8
l8jhGY0/tOgwu2q2N8Onx7wfN/bPgynr74EA844U2DIILQNzSgGEL8vgLaNnDFVeYMqb8SIbuEMF
UEUe2KbKUFkGb9xq9dw7YKfiNIVy/wFUVfFHRDGCe1e4NB6Tar+1k27dMXzimvhcWN2+OmKrtA0Z
hLGdGha2lmKVVlcvXvqzqKyr0DO5NzoQpvkQt0Z5EKyUEX+rA4kW67t+P7Te+sItJVFRok+xOWtf
I/YYgOmS+50aIgVzolaNYtLHcITno45WwrYy3l6aHJpKsDaz1pHkGS7deOIEecs/UARM6LF85Ovk
9KKS3Z5/Jh1na4+l22aXKrswYYB0995B4t9HIZ7p68vudoYYUQrhvzze7Hruy0t/YIFsT3b7/mKf
mmfzz6ubVEVc6gbb/oZWh81/p9oThXVT7oojLkdZIeu5TVcitWS93Il75EO+7mOCbwKqCfHdbWDl
+1r1w1TVmb+6REov5oycChAuQvu2MhaAkTqwmmO0D7ap7RJf9jqSZxQRudvfa+e6SFlhzl4to8Om
yrNefZy77fF2GamxsaJbyY9+tE1ebdCSsqgHe46/eQ3PbbNUwkTXgBRzQi6ezW5fOu3i66wEiaxD
4lEyJUMxQwFKjwjSAXU7HAF7iF85bV41RGTozf1Nb5XqXb+fScHmh9PDRbhcIZkqYUK1et9pvHqq
drDS/DqdTGy656IHfP5TvzHo/Pb8nqfsCmSEKi3Zl2m7Ls04asmNqnK474Zu+OlLzQ+l12zeWTNJ
i7dcmOr3lZNg6gMa4hN00iivzHPZvmpPEIllkrgBJtwPmdrAg701d6ZpB4y5eCZzZaPHHaSdqhP8
KLXpT6fMX+5wOOXwvbC1pUW4ebnIe1mPaJtbm56rgTKqbY5b8BVLdYxn0C+jqTARFiyE0304XxAL
O0WsIE14GD1WvMb02SxlDoCCHhJM9jD5hec4Y08pUJR1khdhQluMkIMTxTdL6J+7lSaFuCaTeqfa
ZwJxJBcBh3+ElnTpk9HJ6FNk3OXf9J6FUP7HI8X/BNpkCk+qK8T0uPimfvqRKac41curTWcNckIL
tWdNhIz9oHwxsDN5w2IPAvTHi830AS/m5ou/AIhXXUUiifdgUeZWoVX0ICETZizRqUcwnj4R3nVZ
08XTS84It7MvpKhECJYgS64S113f/zd8So0VrQKUNNRKC4TihLuI2YnXRGSmGV1jWJ0ehRnjpALo
3k3O0oOQOyu/z6JEoJDEk8wxu+t1IYh8YRcxmhjW2BoH7hXyGwMccAHKU0xWP+V6wg/PE2Ss0ChT
Sv5nThmOJjnGrZcw2ZZsB7PCQwRnsDg+v+BiZ9IyHmoJM+DOeiuZpJQaIcrYqN7sE6uINGe8QeeJ
XsZT+bLSnLUzBV+X7ueO11rdtHrR2RQbNjQamCG2IXAHaq7/H5V+SnB9DI/9nhPivnG/0jsWfKhl
hEt2XodTjUp6Op1w/JbWPQ3jiLvazWku3xKtVstLMII2Ee2WMmli4Qeq+fgVoQKsKj16HeWkhA4N
dlp592n36XAIyKIGM9VIKmhgJOBq49NvVIOr2nTgVf/Un6ZyHvp5P1iEOBahZG5rUaYozMeJcAE2
x4FK16b0JvHuHKZfNoE/Bxe+WvPOJDlL6vUyup37B3JfCcC6jfSik2QKZ/UpgirX0U5KstsLuQm3
3v9o5W53qP17jPq8Dh60f0pGvJepKYaf1H5PjLqKndf49E7X51O2O68/MSIMIJq9k+sWbTeXoxMz
p3ieN8qUgPYgqL20MnB0Mcf0aQprnSj/gVG/7+N4aSzXrQ+ArYNAg8jC4pmAze8JHxzzD6jZFOsV
JrGYtiI78KQuY0Xjc0XjPahv7rppt8mMq3lnT5g/1BRSWsVOzetoYiDKO8MyOqhZRmEFeUJ3YNZY
pJU4srgDP/glUd5QfGwedB7XW7xSdVz44dVzVOY0Ryf7EVBtcYYP3qQX22o82cdLp3gTmOzaqUBo
tznV2d8ZSW7uAFkCGzNuxvNTfgTFdGNJrIa2VPKny/0xrBxDxAG+yYjg+jigNVhQA/CM9np1nTKr
5TaxdBZX5vzKqgLV1Pom6li1GXrhAiqui2uB5C+culPbEC377a3JQi784HsOoXcJcrm+Fdl+PGe3
ViuJs6KB9m0zMhBUjLOk9LIJRPWORddYQkHfb1zg2JJ+hdwVpGExuwdchvPXRp66bxSB9Cs3gEou
8/1w85msVaMs+3/S365tLdYi3mUfGv3ScAm83PJDiVuoTsf+Bu1J514iRH/vGEmXYlq6+95Jbw1J
rn4Kf49kjJZjYZwMNgCgb/eUpjOhkz8RP55Kelcbgp24QFt6+SxwsElshwBhrXzRpOyKXvtyHHOx
Szgo7quFWZK2RfD5Y23JH+IfXcns9AcCjwLOGALX8+XX9uniOdnv2zhk9W08zj/7giD5KCNyS23I
w5E8XPFRGPE+JiRDfIreT2p6MOQJkUzUSdL2152pgW0iX4LW3i5qoFFwxAwCFX2DTBkG6+k7CG72
j09YEnwOzR7LRMHwm3JBVzoOhWaYCb05YOsUJACRPcghx4WOLHJLoeZihwTQgeqJ7U5hjT2vwAT6
1TO0JLoPmjPIvL+HkZEaH03qMQS42dcksMx+ExlVNgqJ9+rOIKuIJGy/nF7L4ZlK+Nkd+hmIdLIf
TxT4CDxYEKTWyK3IGz0qK0yDuEhxMaUjPlV25GWA09tbWoEnY+U9/T9jSFzCva1xzYgv1cGqNcAB
y8q0hKVMtNQQy/bEaoQ/V6zL3yljAXfwqM5vm53NtTszMnm/xJtk/Q8Xfg9yHEHmOGhb/+pkZSbb
AXNVE7kd6JEHQRm8+bB/ZxoaTAh4vqr7DgxqmpEWbKxQWR1eJF+n2zbTqpNmtg6gf3l/q/B+WR3y
aqa5nY43TSP5Pw0ftto2NWORE5GbMH02opnButl3+tHKJORyzgXux8LYAbL0//jAg/GO3v75+Pu/
e00YjSpc/UsQmdgCzTagNdq7S/st/4ym5LBPthPBjBZaAEnhr2xA740lxz3/j6sw1arHuuDlkNIk
O3GYLKuzgYmSNegMYYU3LHOxk0i3L8v7dRg+PBsGAk0GvMwKPAiLV49sZYyhzrnT5VcmHWoYkUf6
olT66InQxciCgooZXWDziq1MtnCKnzU4M6WZ07mv6rFikzmVIczp02+AHbqIxYUnn389kyAH5N9S
rUxGfksa7u5loABPOzZQn1+w21K4MA3ilGzpBOWHKGeRn5Sj2ummC71hFdrGX+XqD+/BJSmAhGqV
7rJWYhdZeWRljMmDo76CL22OQ/+HRhvl752+nmFgZGeQX0DSSZ8H3nnR1EXTeTXNb7Hjqyvxv+Jm
7JfqsXzQELxFHOsO4vb31lXOjej9tFcplPwXVMFCyDqjcWC0R+3aN2QgO8YA86lVmQ+N32YD1gOY
Hfc0iJ07ZJ7TEI8X1SLEjI3v+2Er6zDS/rQifPCOFYVE5fh8NOI9DujcYt5aKcBht67oHRtcXtLk
AOJ5Bh5X8j+/6+UMzr2IxdFvpAzHKliw3c7GCjj3ZlBKsKA7DGnO0R3D7KvVBI5eJKt9KAU2Hb8U
l3BUDzqZfeuTPcbZHZ4Oli1kwXSD/xs4tFRmaOVmhZ6onDSrDCHNCzYyFAktT7a3uuwvN3HXvqNF
nNnFroX2LBsrtat5Z9QRhBY2oHcWDC6Sy1n2iuAOP5FUWuRlUESUGwys1sM92xK3c1WvsvYqz1PJ
WAM9gIQGw8MapdEw2gqRnnJSzLq41ZqqNcqkcrKvkSGGXnL/Ltj/NS/Cd0x/b1xAP+vEv9txeTeY
5j/w3JlbtyTAegudX4UEBI4pSllzEu1eio02ygb7MZGHCTWG7wLrmfPANT5oWM7OJbt4GPeaj3GG
puWBSTuuchmMtwvcAanrmnR/e1/oHZJQwPr3yeMG1VnuHFW1cJbE+GDt/FkAM24SSuHhGi4ClCQn
aH+vJ9/CH5/Lk/FBYJdT/l3YtoqqGZkTdaO3u9a2T/qWkuf8Y+gKUbgPYyTTp2SDMVy2u1mF4rkJ
/Aon00+o9wfSZgW3e1nho7HHxoC6lMakwM0J89UyDYVnCARq4W95CzTWUqhhuk0JOUYAK2k7fw+E
LN97vVrnRpOmET2fR3mQ646lFYnq/20FG+DaZPfJeO7bm7QK6VVFOZp8KkSd2BJvCGmoDqnmG/79
5sI6jRW7L4y30y5biKDaqfYNo/5B1GgjfZSNNJK4BF0r8QV++D0nla2/SUkSMVC/a+B6fHif6Qon
R10os2LxFviOqDJ9O5eLlAjFThM7NTXdV+T+eqnA/1GuKe5pJPciii1HeIHQi9MKqYA0O+bej+TU
8iNC7iZIQKlbsIfAb/rNgUse80md+Cr482iO7y1kG3CKGJApzP4K7/l3PxaT9SiF4yP8z/NV6juu
ZIqqXsL9TqrEWmoPp8GrgRPiK3MpCuTzSaFX55fEkOuFoIGXEGEEOExj6pYa55WOKZOgWbgqa0IG
fjPmYfi9j3t55OQ++i6p8o4K8S5I1SevTEZ0/5pMJO7mE+XAgaE3aK5VaAOOiOLg7cMGEFa9fgvl
M12qMdHpZ4TnMUEPZm9gH/k3CZ+dnhM/IUMQ/XqiewtYp6POjDvnx47OhV95Domf5V3cRowrV88/
KqE0g8GZUAXXblDy5mVI+b+oDDtxZhaPGNICGuchLI6ewidpefM3Q/7wb8maP0WyuBQ2qAETB8Cz
PKfwooL4Ndt0dHnFPVFrZZElZ0w8geRWLyDfmF5yXFm6Hpjz5JJOrFFNGPGTZhkKLcRGioF3Z1wA
UTvsjquDd3F/DP3in9L4H8hW7PgXNYgurCzzUFNguV9Mha7k6OFqx3TGIVhXoGUoHj4X5uRed/ts
fFSMTTgemF52ZDKy90MGINGmwoyWyxP5WGGzDyA+Qj3Mj53Evw5mLCM5VjHiGx4jMxlJ6ruDHOM7
z0Yy2FwchxyXY2yZdMpaQkUi1FJTZlA8pBtxr7aVnFP4Qat8MJcFcq7awGdUPZqHEvK9/ALTYbV6
EO7K60tuJbQAQ4cNra/T2jzL7kNQy5g0oRkWwx2WIp2cWOomWK9p7zI8pDMj2XF8TBAb+ZY9DBd3
fTikFsBVTf/4Tz1Uc4y+lLpoHvFCwGLPwnXrQd+WCQTS9/CShRdalEhvS7UqOcfrRT8oo66E7dfv
u+V/Zb+5TvNdiGrt0X6b/yQTklzWt7ruBEN39nI193s2uGOX+c0KOBZ9qqq5Lqv3thcMVawBU7xU
iBrmQu+teu6lsQ9itC1oRRiIyUpGkcFuCx44f0G5tCdObLDiNyRaRe8rmIG49b4QHBCtpOEArI6/
43IloKxKC1PoZksUgznP0ys3pPDqT1X3ptdtQK3CHeCnsyd1eI37fsFC3Fsoj7ZH6i56wvJrAUxV
IA8PvkvPu1F5UXA4u2rXxUrQCEOLpxKBtHD7i3Vt4cJ/PoJnukwFcONlZIxwYplKiLlEslFbO5EB
RI/rhq+La7AQeRVvFyTC5RMk9CtVYnk/qxrskESr7LOtQMDUf90A4Ou9tvABpWofBRVNR9+n6q3j
mYbAPdJN8edCPDHJ8Cpd/J4tDHFLzslTOMv/gyMDKWoKWqRfGomrbsiQl7Qe4AVfMs7Oo9mlkF/8
JQLpsSIGrUUvcAvk8JHB/VLjCV6/nwqe0fWdjmjbym84Qf5FulRkMFSxGylrfFsvPLGTy5erSYxL
h+aOK6qfIvcLWRnb9g+sryWBN7EJ7nxEOTVWb23YNnb3Xt5CcBLG8Yq57k3hfFnohNNPzoJO0QXy
VepnS5lrwmf3cvCPmc09Acc0PQZcljrEbs6xRXMKnsyFm7yWKTXwRBUAS89u3RW5zeUfAdwV0IZw
qvl8vrW/JyV6kiIBLQoqS7Ca5XhCgTumGphzWCkK9i4lCEmiLgjDarjnNzhjunX6uUHT+0O/yL6y
pJmw4AqClspA5VrbZPvgNtQvXVUtak6WwTM0wBQlVxqDB0AxljR0kNXYX6vyjPecyBK5lbf1dNip
1QxlF3EjCYKhe7ePkOFtPZXLJ8pDt6cOvHMkqRkpyxMKOCU1SEsXNr/Sch1AOO0INMvvwWylNt/B
cUtHuOdbh9+Orsiwe684N4kG1zrZZsEK/JfrQKkD8A5kKbz4zizxbUUBQ7F4AKwc0tkxXQTFGK8d
MWOGpBL5Yo+2Xi2r2Z+moOw1stk2bped3pbO5TPeeLzRUtt20myig1JzNnAkONHsWJim6rZJCBl9
DGhSnukkyV3VkTDTAvOArRW390czESNaoj71hBIvPWvNukz1czk0aP1GcyiuoWhS8oMgdqgPstan
EPvEFvqn67uQTcV2BErXSbvGrFesVLrN4hKB7WNdygMBrMEYtl4PERV0urO8EcDgoWBMilu7RWcS
rH/j3LpTQOMejz3pc6nTwBxQfyloLsQtUAcdSd7X3eOnmdkA6pTTdrTgFXLJiIrzr9iMN/PCDUh1
1l4xXTtahdaJWUAWdkq9B+ymx0dlvNu7Uwzikxl8tlKFZSpDqdcVxdrjdOY5mxuz8NO/yR2qbv29
ty7h2cc0+HziimC+HzUZ3qiwvlVaGtXttJzbJ5qynrXrxeHmPygzfoUjAVZJsDK4vZMg094Na6Jj
VU4Iq4+RU8AIR3nfoKppoGUcDslhMdhcrt+HBoajPbcsQ8lcmBHSZFGL3dDRWaUB/fV/PFYDDJVz
EOCMyM08UknFFdg27ovecsp04m35btMX/UeHVgsV891UDddUTRhRCpd2UhNl2LYTrlUv9zEckRSu
c45PtvBodk4rsuKYiUUXMyIyyRF9QUtvXENKy4mvAOX+gEHi+IRdDteIDSvUhyf4zLWp7J6dgik7
R5p7AMfX9kIibGz6AuD3358hKbE/5OWwrqZW4Jw6J8qX67/E7XWwhjUfXD8KejzcsV4DLwIWeVfx
gAJU5POcDCynh1XJNf8/0+/ud45f7mITHDCO4F6EiE9WLBmwVSBPBLuQXGCRCfCPqID/ZWUBm7GK
xQrn5WTIb2dNmXXyCZHi+4ljKOzJ+zT9wtm06piNoT0AC3CJ5acdpzeaaAVfBNxTRV7p8gqzLKzM
5KTrPIpeFNRKsVdd+M/QFDKBHafgVsxqPC2otIxe5Y9wz5GOkFML5zcUJo3CcW/sO1tETxQmFj3t
mLyw8i0woNUqtcqgr+mZDdaUW2pOfdgMtjQId/PQCYhbH6g0mzMBDAFhLuxpIyRQwxiuDx0FnZku
AnqAzk71SZUDredJ5rvzY6K1a1DqkU2nIhfY5f1lpUMjb/eOQ9LhtdQG7ePvNuV7GejsSR5BAFQl
RVfXWexZKu/KITwC54s2Yrw4FRZwUk+aEPGuaP1yLXyBAPowdIHYot6Ksojre2gceqEqohhAd/Ga
tRnCR38mjhHxEvv51N3GKvk80UlIVUb3Iu1okFQbGeImFB4qDFBXXXgUV4XnvWubCQ7Ca2zJpcMS
+JgiuNvDEoC9RXtJ/erkJm2EPpxGflm5US7n5b/fnOhJ56Ipdxz5+AZsCu3wu2AIvS6aIEBgqN04
hiBdnThFm4wzcFmibKYhXArVE4lFsejPhTeTzhuPsxYchkEKajGLu29COKp7vjrIl2AUL+0hHyep
lEmLLY9ERlI5x7knuzfRsxlw5TrJRm7Q2/zvzVZ343s+QOK5hciWTo7hDLgwJT60JtpwELJm2OJk
QD1cFdTWquP0XrQuGmNDxY1oHUrumccLfmWIqaiMknN0zC8UaqY9i3gGbC5GD2IH5QbqmibdMdPu
a1oFsY5oBwV8S5FhsIaEgHT64SmzF7/LPIygrOdm2WDyCP7V8QR8ti8JixLfFlWbt7Ub9xTVtqn6
cUreP1yMDx4ugzfS9ph2ACamp2MtYM3LnFtM+z4Vf34+9IXl4qKyXboty1zZ5MsXZ3dWBE4D/Oi9
xzfX2ZD7WlGmp0efXPQZbD+TkystIcFwHcIrvniBI1JjYkPKpjdRLoamI1ubTepccvMMwX3klkm0
nrWme9+kyzgeShj3SFzeVkjefUzuBrMhTxaCSv9XT/9YhxvM51V7lCOTCM5lAohFt3pf0+pFriN2
P32l4f+0CIbd1oO36e87Qw7uWmLJu9Y554LLAYyZggdrZsWGZjEb3pOa1VDZn9s/AUoDxiI9l8M6
zGuxE3WCs8HyKu58ar/PaaCnRf+e9p9jjqRinDGAR5/1tm8Awt8lPp2CztRzk3+qIzihSSTXorYL
G3+AJK0twvHSd9g/itVVW/wsuZ1aEsg0+S2QttoYRuAe0VgFGFI/FozGSvjfARUEtbxOhb5em/X3
vY4HNfL7XsyDdUAFd7uJ56MqJ+M+D3HyywYoM/9wb5i2Su0Z386lguhjVY3Uqe6dT+qaT5Rodcr/
7hIBLsiUEzJ9ZGMZsKhczHPPSQEYIDg/d943D6cphV33Qfc9tZoGEAcFaDXvHbsfoJMovSIlmvuB
hMBJaEgcN2kIvJjoVLWzwmLDGzvKR5D9UAK/nZT6cEKWZRUe4pu3afWISuQYQfqFBjgwiZOK+8yk
avr6ZgaDci4HGlOwPfIVpns7TH7D4IgPM9aNQheSE9IfnSsWdreekXCXrEBdmnSacUJurrrO/ZDL
mrfmyB0/LzPuqgQ+J+ANp+2lXRvwMfNs2JUNlBSoSaT3TC5TbN1o40D4CNN5xLg9upEHuk/FCetg
/6kvxroiR84qXeR52HDV3TCQ0hcwxihY9e+jHfTENv08DMFL3zd9b9+5sg/WpoVvVZC3Jrp7FnM3
iA5XPen4Dc5eyNJE/pxLTaLnu9yBFocGRfVderGyFBlvu3DUl0whlaHpWecL2U79dm40S4FTBz3e
q55Y6Xz9VMpj5ztkm7pvXfwJaMDWWUeK5vDqZ2wWdGBk2fIRn3Bm1KRhmYRKx4itt7P2mA4qyta4
72YwPvilWdkM41IwUByqBbEylR39b0DUdgsqteKmG+osdaHqoKRpk9DvElDxn+gEwix6ejz4Lb16
EcKuPrYvvqA/PsNTrbUbKsE2h+mnDFxQmMpfNHLI+FYE0qfTSWDdLRle7eyPEdUyxzm9d9ArN9jT
D1j7IhaBJlqLl5Z1idi9/XwLZ20buPe7x1QEJCHDpoNa8Kab9fF369E757pSkmvTTOoLfTYZS9X+
p+CWwESKlSqOCLZhui1dLCnES7A6KDKL+8ipXuMBAe+KUn+EnvB9Bsh+M+CgJH6h1lfgFn3eCCzh
aAvCIpqizkX63n5e2eClcgJvqIk5xtFWE80tcJQpCrP39WVbYV1f9vVfh2Y87RVpYUfpI2nbi988
I8SwKrbf/xyXLcMiwVqAWxgj4cfVvIN42aV1+Kt2LHmGroajE2JIeUJyyCjEXWPrWKwNiynpbMhm
xn+RyvuoOXFkKnrAjIxcvCldLdySGyFV/XQSNv9RDohgdoX4Y0KE8tGTFdwnh7EAan61+R4aOaeR
KFHogFJtJT0Pxp63j5l26AkCOqWA4Bp9xtLUz4LsF723O4Jhgoxsk8XDNwir7wtfJYHa8IC2ThnI
lw8gmq//8lxIMxEcaEA8jsyOn50tQqmEx3l3o4cxtYICj661zOZ6j3yOJ5sTBNvTmMIdMaDUIVla
3yIGkJ/C/osDmce39efWRXMKP0h/dvVz6qmUNl3vzVmMZCocNEiYdLkEyMCdsEDGn+kODQZMqoe2
/coreIuEmVu9eV+ES42AkfrH2464SWtLE7SkHFgrBhEqiEtZ5S65evzCXKFjEfJRVpLOJmxe+0Js
Q2HWAaNhtmZImnHWdtp1313sKMCl+PIwfYRjV7AKyBZvXvqIWQJdEG7gNzOYP8B3THHx6cvTg1/9
wU1CT8/EU7U43IsIUs67wo4MBuMveyu6nGueh9B2GULu3r9fDYQxhTTRiWbP3Pr65ViO6s+++zjR
3538GqSy3QAZIrAc1UdDokO0G87UfBML68HvWU0kdiYyDNdLWDx3WYbVR5KE9iehXUE0F0rdM8TA
9LPMf4r3BbFZnPTflGGPsch2PRxdIilXqskfjkA49XsEfc8Av/FNAs12ggef+/R6kaLRBxkEaIqe
2KSWXZLX0uWmaMXVqdSxf9VIbIIZZ1iyyWzLYTUfls3kDk3GQXlAOH92LcwI77itSZMNiTzqQGkG
AqRm57ylpq1E9zE042mgQEGnQTapBZPMGshoCF9wdyaj17YzP5femDRMyTP2N8nMqZ3g0oL/Sbqm
KTIjhlqj3Hl9ojRT6dAPZKrVfQW/ungRNJCt9qHZqIzbWIFZGCIuG4QpDMadC6ttIRILhWZyvd/f
QtO0f/kFPS1lw8TJGjghOGqRu2SQZFyBks4JiKopQLs4zKl8s5MpHF4I//X/Y2e8LHgESBl2Lmyb
ARFIdwXTKiPTjDG1zdqBzTczlq7QrcxAe6DcL44DUsdim6Lr4SP4MXZHe52T8wdloLTYZF/2u5ky
0uQ+z0uMCshqcxaMiwvPLrDWPKz2U/HpRWeMyYU3yoEulR/zHw3b3FGdIboX/9HbnUZR6DzG0Zef
yFFucJEnka/AupevQN3mNED7VLzpLcB61HcjzJluZZMhzfFvfjB//EBPcxv26wIs0rWChurxFFSp
Y6/ams95ozor+en5mmeQm0v2YXrj+jS1wg88GSzfeql8r/64eGGncVDBR7OL2hYOSRgeaKlFnLry
HyiLLW4rbsIaTE1O5x6E9NM+aXVMqVxxz1uCWvUufk97j0zVfQCgWXWqyJlJpaMtA4bJiY7FAmMm
zu76I6AmiG8bahcMOR/wLrYNI/IltLmDlAAissa3rRUZXLqlCCkp+uIhx5rZn60I1wKkUguIOlb7
28mLeBNtZzl7MaO+oVvC75QZNCYRbj9NelGTrsyIKPCy6YdG0McmOz+N2rYbtrllUiB1Nb3Cit3v
/XOvGAnxdDKgsYNq2zfscIFN4fSYke2xoPzKBEK9fXUsgj54jf0bCCH6c/sRBC8BE6NDyNoC3eEJ
T7Yf10V7yPzfjuNsyskdkr9NO0PYfj5/JB7XvdE4YCTfIlCFtLw1MN5bNZ46B4e6qSnS4hrIcPS9
Jf7PHbUmxaa22slTPSWtw5C6L75MuiVhkzwaNY5GlSd0D1F23rvSrAOMAu299ari68K8Vdt4Cgfe
0IMgjLDyTR9DcRNJYO3HXmf1UjhHPTZER7kpwiPU2Xd2SIAX1dG/5on48IwFvkytSJ/BoXsu2+E5
kNQmbaFCRdX90wn53vgqTdKxo88Owaq6LUnH8sJr9lRV+wnkwgMPu7ivvJSTjDb43wRXzfmLyHcc
o8eQ9jSxJQ+thqbmsisTWkz0IupqPeGt+cnkDqV3pmL9ypgwq77ckCHX5/nKGDTVlacVFLVGE1SK
dw39rJpDxIPo9xpezFWmrtPVlBjGKJJ8DEhxu39aJBgC5+aEB882IKGRmQJkcqM6otf8pK9vxpAa
X7QTINbklk+eMHlXL1lYtX0gXZMsWUIPrxPOIoPpv7WiRTvwuKA4CbydQdrZ+1SzpNMDy8tQgkdh
bhOQDMl+dy4UXOtQqZcu7r8rc03uo9NOO/ttwWBemmp04YkD7dAitjxsmMo9U85k0tymjBSHWrWD
Yh92PV1Md9bOEi/txs9vcYfaFGSP4s0JN7L4kjO2CmLDK/ceIh7ASnbGOB6qtNL7xlFvMrr6XY3H
cfoUE7WleH0WKN+q27zVNzDGepzMnRq2iQi4Te2j0zwMQzuL4Qu2R84cCOT+3K8IEciMlQtZqOWj
lmdKngudDadk8YIrffkl5qp38Tg2jRAdkza1bh5lq4OeTNeSwSCPmKKI0nH8oRmIDbJQPtt4ddJd
bMJrGx5D9iBRN1+VWT81lbc6iiiijn5veAH542H7ec6QDOdrzCNfLZ3vTSNan79ettBTHrb8ieYt
dvT7lWhNcFde66YYbqN4lqsOvBpqdpWO/tKZGWXA/1E+cPwfnplNp9772KcpQafe13zCnXdWw+ql
rbNasU5awrBliSbMqBTspJMU1QugtwR+IUOascKo0hz+g/BSK7LfJgQcnZHt3HPEMevVz6A19Nfc
fSYGKK6NsYnDUefma7iZHt11LL76RfC9x804aePTfHK5pI/rTH3b7JdAlkyRUsp8HCdK8sTrEJK4
MMK8Lfdx7IEgfwBktmiBboBqUMYsPGxmx8qJlSgpcNhAQy6l/W/Ugqc+D/63uIC020jcHV0gjhn7
YETqLhUNpKyBe+81XvM1ha+llGLFiL7HmZNqsxBKiyVkVOpIAc1IzgouqfrD/HX1m5dr9ZS2JbKo
l0xpgVVKFH8y2MOUUCO4HZokuA9iunETExrIiGEW0IMQ9S1+znW5WUkX9zFypsGIU3cr6hmO9Uzd
TuGJvuMWsqmqhYYTmVVOiYiNszJ9cFRn8ntlvdlPWLzO5wTIWb+ZDwEj/brvJK/otfswLkfa4pME
7z5An0CexdENzL79rMfN4tz7mAGeNSAa5bWmnFnwsCwN6SLZ7lrJ02XzWokifzJj4tbL/4vOpnKA
uvJViGGaWsz1yqTTO4UOlNdrNxKZG65E06zl3wvjRZIn7VPR3FhkRFe826UU/HfZKkO8o8tUeoNz
l1thGFmQIFfowdZEcTmlrG6kWPvdey+hpLkWoZeQrFUWsE1uu6KgJ57MLEHsxbpyOYRyaDphdLOB
5/VRS2ZYkylAlkjsi1M3kNxC79VWJrSeKtYheZxDtCzx2UB1SAdyJetqDUmMLKmkgEN9J/f9oPa7
9iY4se2G+XwMV2l4uE4G6WR91bPde/YaY14Fe1cEBRTkYWdYRT7JwaASAgONMlycoay0Eo6CsM6u
w6IlL1dBaJgGanZC5mcmoNS7VJzxWXXs8bFiJc+7qo0dli3+kYvgHuBcTLpzNhtNbwiW5W2sOPZe
fUh7qz3TFNRY1dFJnYla8Z9tGQiYfhAmE21B/p65nGhNQxpzjJS1w75YbBQoDODN+OZrpaZbuWkL
7/nifWfSlh086Ya8lFFbfLe40+fi1U21tjP+PMWfTRrJTYLaH4uigDu3/nB+QY7ZaxYoYPnt+3Dr
fAsHODpqF4E/o5E7a9SEkWm1HVDAtKiT8rfExWg76OJbjeRlFTGA3clN14Wx+lsoYJut93V/VBZo
kqaUPtq+tMFq+a+JPkuEwtESq/QJO9bujZas+jxjcEzVDbnzn7xtU2K8l5SwDzB+vz2wFnXqPZAF
Ww2DiWvrlkPgLzBTHADpYlniBLzf1FqxMMWAYIUzQFNuIGYCMGM7nJBX8m2k4crBO5QFFRgq84Rf
Rsr34eBT6UBH7ygn2G+MsdqMV9K9EedYqO7mN5rxXn27PSGQsYLZrT9Zo0mE4GpMd2dvD8lnDnzp
yz/b8QQCBCDux4a/YyiF+KKDQlsNcC0FS6T4B41i6pRxO8FPcgkveuNIpVS5VFN0b27q0bji0ZY3
oK9y0qak0IztgW6NQTbqnA2ZOsWAd/NALCfIWSZ5gvR7Qhfm68f61j0ofC/Crhr2nPZqRiIwId1A
m0QOLjqX1EkO2HO4cgvmp3HiXv3z1PzI9HBQxHTGnI9OqVw4JYo3XCifpkHQtGFb10iel4aBhKDP
QmRzltCtluqDVNbCBOJbKDbKuMPLCtdh26F2AX2Aq+bc9YnZCECRFImLZPk8Q7axGnAprJZJL7SV
GVdIVjsrz0j4R3x8Rs5g6ruZSsBg57rZIBvBXte7/XC/kf0Ctf1sGwHiFhqDU/5E8SfYC683EDvS
vFENKa8ux/UiJVEHEvJhxlZb6ZfwjF4tM7czydRnlvzfHiZXEtqPBg3Ncg4EIvdiU/DX41UPfsUE
JAe69hUmwz2IjH+oKm7SG+mwnI3l32JHWIueLKFXoZ54mc+qERVfYlwcNqWh7qme59MFawPjkfcz
6sb1LHADGZnV+jc6ErWIREGpNBAycvT7y/17nMwL1UDaytm/zFrEd9Hk7K6XLujZQDnAuZ/BycnQ
gEu46zawL/7WTmts/1nruJp0G11e9LDGmEgCxccK4uo2BkvZIDNK+Z+r33IntwU9AAMGQIaWBQdd
lIacyswsGLaaqNNtuaF/8t/Q9p9ks/jxFDorWQ85g7Agfg3FgcCpXXDj+pRHwES10v7URRlkCQet
rpfr9/hTHzSDbzz5T3i7VVqucJvUiuid7sxuFj3so5AX4JGt58Vb8ePFrD3hbRbSwZfj72VVEmDS
vCKuNBnAXtkrHPKVVtb0H5OQkI/LwmN/4pTrEubhxh1SE0Trz6oNavwUWLo0zBGrDoV28Q8uXS9Q
kAdO61N+ZHRXhVbqxbx08ga1XsfKbiSSda6oAr/qKMsG8rxnz7WOMfH5n2yJ/Ngn8cgtJYaAYilT
w6leosnVkRoYX1Zw/BL05fUu12PKWBr1pqwuEK70KuFExQT0R8kNyi7D8w1+lFRysJCXvOFq2Vv4
Z2WFMfFpE4uYzO4mW3YKYTZFAQcDRk0pzIgoQecAwzmeqYL6ASVT0dhEAOJuqucsx4lc+OPchMx5
/OfI+2kJAFqt08oALtpOV8RvU/4dCwVZFStwc4XOkmUAvSIgpcAj8J7VciKbliyZnZB2gJzk409G
qELGdAhBwIqx4JKmmajxiDNOcAflr1/O4LNIsRz8Tc3BG91Bi3Oww/6pKdnewE5gfX0ZMrDX+L39
3oGqo6Sq4cU2Se78D8AWtK8X7DPn1qIjyOg9ZGvAxiawWK0HMjQPEGEyNqQjH/sjB+6wRp4n6Svx
JBIMQoWuZvGA1cQBmWYfKkM/+GSL/qUBIAPXLKr6NmlwU8lI4HoT1BZLmpt2EEZEruAIuXhojN2f
BbueLpvS0NfEvhNA58U9jsoT3mF1VvxH7WB7B6ZCD+ZjShKgSXHWF9CKtAdZQszAYh/NNKC8ouz2
1V5cKiFghHxPIvWd1hxQNaTwoKHyWGfYo5am+8zQjZSmL30KogbsGxMogxaQLR3xfhUEuoKT++m4
+zysuX5jBEB84zBqlpzJUXAp9+WTIHvdjLeZZ+xTD5LzbVoQJwQnislcZnl+7tJiSqHZph2XHqXT
N0rX91V/kYGCkFn8EfhuXtikYqW19QyYhDmIlCXso0DbM0CzHVXWKYhpZS8RbYIsnBWoT0v9Z6RK
Hxgah/qF/WnQpbJWdHeTQYzq652v4UCkVA7sUX4dg6Mw33BILRWUTNZE6sYuTR5JzW/bg811Ed6N
ndRJBy3jDYxlhSWScWB8uypTZffI3WI4CY+Bv625Yvata09bATtHF1VotBI5Q6sWQ1ZEcvSKQbP4
rwKVrWQLh4bkjxvW8lgNFq/gqxZXQ59ayQUiWGbs/HEM5NORxm4zs8sQN5us1ybO3mLV/JwIZ79k
gGSS/qFAtkmj8uIz7LpU1B+16ZWFrYG4MK2h0ULHYnY5Mi539ttSFgzIgBZkgY+unag4K5pFEDQv
mQtuF4slsES7Ds7Ss4mYf3XXr6FhQm+uo+w6y1737hA78TxsMKbsESCHWzWe2E3QnnFqVi6IA5bp
15HHj80pOUJarBO7+m8fi/i7+hO9jT15Cqk4HlOxGuVit+wqS8ppPNFiPsg8zp6ysRhykoIwBIX6
3VisnBqFiAVTBYp1lt2JxAVslyxc6/mSakmPJfhb9qCTWzBWwjpYTJfEs3kURzOYdApjZoKWIjuF
M1k6Rl6eSJ1DzS55oXKe43OY+71jZ1en9Mbg+gC6YpbqFMqwZz/Y4+7BneKb8KNXAll5bCUriE3z
BXRDXKy3gvk7V9g1OS5sttWimgwJIYb2uUtsn5Frgx1T7nY24BMQMjy2Qo/NJ6JPi51Cwshu5ZFD
EG3xwVP+tllaaJJrMgNCj/yOZ79Pk5MWzaJnkmfgZr4qnQZqThCxLoYWfL7c5ZbiEmOB7gocsKvF
Cicb+EaPGBoS0Hql8XxHMYOIDjp6qApGzVw7WXyf9WIndEWRrEyAXJD33X0ilo4E5pE5YS3BkGfI
ND7Ccs4jBnaxhjpsvVW9HjcLepbvRh473mx9riVOWrbX53HxvBIuF7fHpjaiZl0AvGWN6Jz7tBhl
T2d3iaW+vDJNdRjrrgm/eviQhfGgvF+ASa78YfjJij83JuPSgJo+iKm+yBovleHfajDh4YRfpRnp
is7/P8cjpALPBVCt4uKlpAJEq6/U5d9JBi+KCDLI1mMg5+bhfoSc+cdGo6VWVyKIpISRZwzrCUH2
MTKT3HgXz+tBme0yTwGG6keglMF45eCdsl8jmNrJmVrGjdNikJ8WSCIa3HGW/RbfnLtCIQptNtd2
IWIYMBbDCn1tlGa4rDZfdOIwGY1nPCwPRs1dWmq6uEWxxmBads4c7FjZ32agNGn7L8pwcp+YCVmT
EOVR+BjBWCYeKo1QzqUvmhTObp9KO9zDum1ov4PHDbZDsLE9xGaaDCgNlZEMgqkEdikCndp5M5BV
j++9HEOeeu0EwxR6vg4GYG43OUceHFy30HbEeRGJrQvhWDlKHTMkuUK6TQijV11wMbShhbkXrvD0
vDJyi1YtM+Astp1JRf1ZvFp/aw+Jb3+r50F+13vtPMxczUZrdNYC80QOIripV1L4DtKZEiBA84xY
+wx5D5gydmUjigb2GmLm3CPzv32Qbh+sqE5Fxk89KvNMoQANzMFXWwwxU2WeMVHQawqmphksue/J
lTzb3Pe5FjMtRCOwWkH/KFuCY29Fili76jXeiSbMQTZcSpXVuHxbkk38+U4pWIjTye76q3ojJukD
sWr5mWlQOIu92elFqGbLrjx6fL4bngg2ygYlvUq4ORUN9OoA4ptRQ3Z2X0K7LoR7vIgs7OX6sUVm
bvjJsKTLdoFCB+uiPWGjbgv3ncp0/+c65BGWF2Y3KjqoiHnOBySZoKZ1MmIq6X6vQftErICoUlwk
c6gKtVRsQ6O9ByW5Hy/15177e1GKiVjVEZUiOjPTyP4AdSp/2YswedfUoWIoFo37aL89/bvoDAgC
eOenHVpdfDP/hCFVac3DGm9IgA+ll6xCMd2BXxCj6Wd3Iw9XM3prqx3sMU/CjOowaeUWepIt50Ja
wwQHyBnE3EbHIGnXXs9T/vMhZnrq/vrEmUtJT5Cgy8D39tbsaO1qqkfgPX7U++In0DSnZ1989sF0
VnTWT1+fyG1xsOwivfz03Mp+Jif8JCLtiKum60f/nO9jiVZpM9rU9Cxd6N+6MmrEzYomZgLzojhJ
EGJV8JqVRQvfLNq4c9wTpXfOHPAXYp/cP+USMGwKd2/BTMpq9Xh6/wnxmux9v2a1+vZcbqI6EJA6
0n1t4WLGc79sLEC7p4BS0y+VrK0D4+FSrLJ3nAPCWz0wrfzsG4Pg0Pvmqyu6/eae+N1RXaat2ZK6
jBAS4uQdeOo7uAgw1p3LiRHUnUrZAvr2y9VKAakH04EuK+WsoHtmXTMVZplxyNPDKZSGpwAkW3Zd
02KtlcXv35w6VWjp0Ys+kFhnrCwgGl3TU0DSxNwD/Y6x6gddhIqESjhcpCN56Q+dHScKZAJ+D16K
yNv/CPIxe9GSllj8KkAj44L4EmXjUwQc9Ruc30g06HE8vVDnclca/bOHb+SEj2TBjtf65vci13IW
8prEze58E9D6gEm6TrmPcM+JMx0SQjiMw84IR4VCYp96NPr7gVxnvwz4tc0b0aJ+RYPZ6+dysNCA
xgPL3ZzGWRfwff1ivEYC99jWmY2vJbBj8YifnZiSDHwjIqJWXEKut3FcD+cwLvtOegljij8k22R8
xf+LS+4j+hKYfbLekoHmlgJhrb9VkYdCaPjA3qkvBJ7hakr2Bqq3IGUyy14KGolU999Bh2orr4h+
1tx08FukHqPcr0s58tTRv8nz0G4PcyCn/2SzSCe6+zctD20PdYOpQAEvRV+x/0cJHv9OIwGon0/4
KoCj/ZpEDBPvGMAMKIDdbtGsW4qijvt9Q+maAlgbI+zM7gDnymuEPusvX5kJAgSCBZJVVqLELCLl
kVxF3jbSn+ZO/c4V9SbCpeiPIfUH1C4Z6phGOxYcO37gRBbFmlLxufV2Q1FTlzcgZCi0CAgpm0ur
vcWChgU9jd9OR2hFc0ms20gz0GKiAFxTGACW30947J6zZt+OhK3kv5bkuLVXJQ5btKSnECtUbJ+M
quwQWk+HYqjsjcGAcH9t6mWludfdVSUDgaCDrhYVX6Mb9JO39h5VHs8Puh/OBsdbNlJ5+sHAHcA4
8qA4ICVnl13bflbMsfk+iTtz3yr0ifzNzZ/cWDHh/WFNuDoadpnwxYo0kfOF16QWOOB2KvvN8x8i
5zq6S0PYN7TVUWjHFek0f+apA7995Vkj/9JbOjUCh1jXQAdTNnHLEczgRChfptA4Qv89DER69UY2
PTSVMFpf3xaaXkEGBnFFH7djkNjbC2br2QGAJWnHPE8NwHray67soLmx8govloJIWzZgDXwpaPsH
znec6TCDDKeSVuCByuAqJN+HKA/Zs3HPU/OskvT83S0pqspv9YvCGrcEFyBclVQL/RFNR0YPQ8hT
IINQBRBwknO2/YD1LnM0YjzFJdS4m8muZMzVKV3fDmmQkXp3EvMrQMfDqZyW+oDJWRV2Vm3G6mJM
D4Qk3ky1zR0xkl1eqxsi3SSXnQYEthyTszf20H7XFSSmPqnI7pV+vxH9nxf/xDUMiEgB0/lS/2Ec
5n5w7EBtgOSOj9LwSSExbrJMyjr6vGVDYP1HUkCShWMy+Wi7EdRvPEosLqGaF+ss2zXmBaGIpmjR
ooov4PJ7mf3Uf/dB6vHm8PRykGevEHb5XEBmnNz/jDpe3nhihdCnZgQG99Twil0aOtijtc4cw9nb
katMbmSgejMSD47W13XsQOGEJ/f177QFmVywQ4c3+tgJa7LrPn50T64cd/3O5lBWITdNf13YC95I
hBTLRJ+mSZGEVjKv24kJhLl72yeqyJPnkuk0OmB82S8tqBRftJRON/4JBwYOQy7Dfssywa85p+2q
XrLIl1Bz12A+SEJzBj1igwAkWNM2PLWI5tFPIOUPgWuNcJ2B8CByAujU6gCchi5qoDGYywX0HOPx
flhgA1V3ZkYv7RCpheKBEHKOIskuWvR7liI323TqVW/t+UOePV4iEkmWEbGr+iRXw0QdB+56HHMv
N4Wj5Qnp6uBqqAO2uTahKngIRNEg5+ZvBMu96HsQTR3g0fVME+wD3DZwbCje6h3rPW2eznWsEPzB
5nm558AOlxGirgf10rLMGc0EY4eRrUiuPt/y3evyyGIA4dQOvth+VEmQaUy5EDj6ZOjBFJAyq3I+
xqO4W4uYEX0VCxD9eN3uvePkJW7DIztJMMzznyuOwc5FC/KReDqyQWMOh1KqqxbbEALf8rIWptu3
2FEUlmWiDW7dXWT1zEY9cKc56/+0wzywD4N/fQgn5421tnSmZRuN45cE3vpujw9wmYRV7aoNb8q9
3nWbV9I7r7qesFx68liiGHB8K83Xi0N/EHsJlGi/VeUQqke2V2mTjXl+8OmB5sPenvEcRV+IEn2d
zQjdrz1cYOtFkpR8BCAMrSgX7NJ/zCCYANoKymBAaILlEHRHfDtRF4pfRzzV+lp1xb2EtP3WWxVJ
XUVHGsNNbFFwxPh022fg8oAKzb2Q/jsHVocJoEn0aLvbNyVHqD/NPyAnPQH0mFYda4aafLdQ+iRk
whOlhuaJy3bz8Nud2wxRQWoW/MflADFTLA4+5gqHnLzLkPr+AYd9QHV4J7MmfzUL5tE4a/RKiKLn
x+IQxvCYs4VpCo2GlK+D4mAsRhoEdtjzAHe+N1/oLhCfAljYpSIjl6Ex07ZWrPqW0uvLB1e3GncL
CauAFf5w5Xr4dOV9/vWU6nt2N3Ty+MjD2ODGctAiyVXug6s/g+F+F77M9fj5Yl9e9ZCNvCOIPq7V
q0zagXEJR1sg3LsJnzSZVjEzhuy3Rl9ti760Z7WFKdLhEjcuiKopHMC605xBib0HiAtDVB1tc+FR
68jS26OClTGr3Raiw8dhq2r01F1QkWaAgaHT/ZlSAotC5kTqHFlw1nrxMjJDhnd0h8iy43bIcFJQ
27jPsUyBzDqCwqG6IpePJKFYwYlq2EXBc1VEQU5qLnsYP/2I67tCLeRUzPaDRus9pmiRbolYBTh1
TT0YRGWQF3WWzR90Zafzu49U2uYE3nzWAqvRIZKXRoaN3ITpOyd3dNh4bET+FGuWzlkiy7cMrZpm
pb/wGwas2ikZJXViC2PauZnXKULuZja6OV4pOH1OlwB16+zQUvkIfEv2s6BpmwhsO/T35EMrBxub
52dUOm8R1KXrQ8b/kl+3A56kTrrVFfM5Ludy8x3KfcLFQPW4pbwTYWHQc3cnvH451HBJgrKXnYo5
5I34o/1SDWOErnIxXwylVg1G9zGBtok6L2YgiAGK4cmtwXIZ3gL/sxmM/kgDRwF31bhCTjaKVK78
wJCGn9RhORsKGAzSYumsBosD+Wk797y+SnmCzEiX+0A5ZI/ldb1NfbdAK6Ukhafx8ZoQXITO1vnM
uIJKPsXOqfYMHejOOaA9lX4998t3leRJZNH6vtSqDZL0OmTQPU8XhnybJZLz/L54T/lMDbPPmLxW
14omgKIrDiWLminfMFbaOJHBApvcipldWl1R5LvxK2lIaehrxqXtHxNLHxiOWPSeCstZ7TZfPJ4Y
6r29xrtD9vjJgI/apJV3Vdolv82NMMqD4R0aVlO/GBhaEbY+OcbSgqfJIctBMm1TXl7mUlEpDq88
alOXxGfEsKn+boSzOTcD+FqDdJCAU7ND/qy46VQs9e7w+jxzI/FGKha2nJe6zVAVklFgeYA3TZcB
ZyeZRQ3yOwHtDBq4mLrKJW2/cMrhvCMxfynymaz1NtE8538UBc2d6BIGIoqJnIq7K/TqC2mMBznZ
6VXGRUI1IBue755hIaHP0PQsgDdQCBJkVDvuYMSx7u05u1DDXqj1tp43AhsJBQoj02avZcvl9Fwp
wDoOVxssUkPxFayDRyzlxIvUDnFZWKRYxh4ZTMJcCbb2ffD8owe0dxa7Xqz3kykRDic1RUrxKQZd
oU1R+zqQpUn0YeZkv82u9+zMTYarVPrVJT1L4w01OBMVVR6nGsZEEJj0B3/O13/6YEz8CemFkouC
G9i0r3W6zOqF3F32IwujSmwk30fA+hYRBUL5ZAX9gS3LYRuOkCw8i+SNSM35klX/dvCcWQAsaxAD
wxCHPpfAt0vu6ekof+YNP3gHqWorCrfln4+kKyo5aL1ICDca+0xKWxP77msBgSk1JLjZF4v7tgnu
/7JY29RFoGTDZ5TCypDdHxUk2fPAwwTEibZp1AYZJTwIbW4eSQ/Mt199cvCM5MoZiDYYZGRXhzO8
G3NoDlLuMnbTe1ic0v/iHerGY1vFBK2eo0uMGiAGEshRUbLRCSKMNDX3avJXVzd2MnFqRLAKqef1
AtDqXDmkpMZT4h4JoYAxANEIgmfbgs9QifaGGzyv7AgSjcq7wiL/vKxq3B6l0MS2yTAdlZPXmVR9
q1t59/V0jTb3tznFfBoG23gq4w5UwMoFtpUdwD94SSSIPivHe9uU5RC8Fd0jO/Fxl04CR5JqryfI
D5tmV7yXeRs3QMA2mlIuV7mW1HD/yMzkv64i/iN5rQyYLnkmc8oPAxTp+tO8hEgu/F2re4bkHo6Z
ZIPATLFjnulbMxBUHSO3c6h+DlIYr55yrJEtr0ZfevIzLkzBTb26Y+H39JW1nKGj5f7zHgyt7Qqn
GlSgrOEGOk/3UUwraKrnLBmjI5PfhJ0sOD26lFW+yKCSdKtQSRZtMYs2Kc0jsPZSx5O7vdwi5w+r
12IGY7atENZlrSwR6JBGETknT357PUfENbo9eNBnJS9+dGdlLrnY0W/zEHJcUIYFHDtQaJoAQqma
rjTMlJ6HCmii0U9ELYaDIxOYArkAoe1u0PvQfRx4qkfLYLFC7b1k6vtAkYYJyNpCEbzgGLKY/49a
MlCrxYPYL1g5loYW+KmDc/JY88ydGn3Ee4A/cLQ4QYeH9JgWU81zTn3UCNb7ELmMPy619l95dIFI
vPVyB3jQJ3vfTmYEromFn1MjxVMdtpVZARNJlFBsMdLnaDW8suS9qKWmAwiShUH23fLtiN6W3cqs
D+aLJAr5PM/zHOFBv2DKSjjWhCaEBYGe0EUo2YoM+s7vy4AK7gSK7dH/h+9ehmBh9V9oqmzhoQxm
JO4Om56gjM5uP6D3l9REOWxck9CwasKKg7H81/tK5hL7D+rscomC/iBBQ7CW5dXKgMhNOkibCxEl
dAMVwu6H5K/ADEbEIGO6IBWN0kjO1obeoK742DaYK2aVPUiuVk8vQPBQ4sGwi2++otUiiatRt5nB
k1B2tIrv3eZdK+8cj+tmkYVJfZMlo7zzF2JefqwwuWU1LFmuN1uPk6uxPkybaFqgYVzzelRR4XgA
FL1hHOyPuLZBrpkvYJvujVoV+35c0VMRKd/fL5DuP7KB4/FvhWdMsQITDwqtYfvnCPDMN7ZPVg7B
cWh5uFEgRMne9c5GyRKcvJOzz2L9e00z815kT4ooEhRkRP2FM7KI9Kz/Mb/l+v6KeyZHUfgQma30
hsBUekum9wL66OEf4OQ+77LKK9Yfg1fQFsw2wkeKf/bFrygzTP09EE25FvLOlLbRN+LhvpxFVX4Z
v1lJyTfRA+bMy7ebiRmLPL8fOTIcN432kzhsx0LDsrlf9ETmYbMBY6Ib5AwajKC+cxEuYHbWUz1c
3ggbR8pmPSBLA/X94rMYpRWzKP5ZkTje82rz5z/dHV/zzH3uwydEoNTLKydMIoD9o8weEaaBtYAa
WA9t2P2wupH+8uG19JyjBO1mpSTogp49+R9ed3Cdc3pD5ne+rDpjwJ+ySnEzcOg2gXF3oHC+3rHP
1wUQ6/zERLH7KikRMvQVnI0u7NMpeERoXd4a/pJ3ik06yo9Gvj7yyTEbU0yYC8X1Tns96b3lY8Wo
W9KQCCXwhYXL345QP4mnOKxb4rHQJu+PXhKejbB50E+oOmoc+opmDKkU1EIWjP8tncpVndoC9M5W
e9uM40ZWbJn1oTHtdno9pSvdzsWZzR6+97SFRCUnwEgLe4ZkP7KZ3reIBAXB/zdVoqAol4IVvGa9
jO0exeboS9bNP9GxP434co4LEqNfb3B0Y6plwiTbS1lMaXaHAZDeGHQ1YX6Z9zHlKe5H/xfHCtNo
ltMSNLxiGjhXd23B0eCIybvbXooOL9xMtFIKGNKB5XpU3H35lRAajXLcPL7ydCrZRrB5iJt/09LT
33TNR6T0XpKojaVHFgqs/efKY2SyU2QMYGcVeRnLMzGdJYZVI01sgsZaR/Welu83jUOiYqLlgENp
lz4Sb10uhtjk7OU/r1GbkSc7UcI+iuE6wGI5wa13UqwP8ylQwI7oy2+zlK16b0Pgt86wydPvFLQD
7ALcyQsh/JC5RNmBpvJe9AUJlGvlCqxT8HZbv8kbbN/jD/h8xp4AkgyA8ZWCI1kiQFuIXNMrzkUT
YR1zXqrBHpUTYtgxgbI0IZZXIf8qsQpSl0grCGs97wNcajs38FIiCdO0SQ5fNFizr+ZVqcsAtg1c
LutuZMHq5kHAF2b4ic82HCyCIVFafXk9biY3P4xLeqdYaEwhMdWduGu0pKk8a/OoUFwvUQVlWAmO
yGRUNE53/GBXIEVwbSAMDZBcsGEwik5Pwpji2LMTPYg7OB3u9KE3CLzhFtgvRUsuNcaR/Baapzec
uDNTqK204fKKt9m9fPPgqWu2hDaPxHyCh/0mth0BQQJGXoxmcN+a270Iea8CBdLZw5WWkHQJtxOr
AFN89mWIzebh8ri0ao/RBqWVBmthCyRktvqejVmAC71jGy9bQf28eCbYXelhdxr9V851sWh+hl+S
NQD42jqIw5upEk7q8pm9qVrM9O/Slvssj5fmMQvt+XiICHVrTadp3s3L26L12aGdCx4LV59JuPvW
qH1N9V9DJnBogNlYJiBtWPZGzZbt98dKAexqh6gJontx65pEMVzb6zLghWDDOkmGqzwpeH5Vnfj+
F3k2fTpovm3FQ0lHcWu36OSOGWJ0ygzWpi59KDpEYnkQnieZE8JeUfoTtKGb8tnwdfJQzGEaz8IS
PIFzBmbUhgrTtzLbvJTzJiNqz90pm1k3up3/4mhx7J9ekgJd2SrIRV/dTu7DBxftXP4+Fd6bn54z
hqQXsFIHQfJ8Q0mJUwsixoRN2RGtPcdhpkd6ObgBIOUX471CMDoMjBHomOFI0XfZvow2k4iet9iL
FpsjqA1mIVbNy+xU5nyMxSTuoZmQ8a/QvzOjhfpvlXtzSS9hEf6hYIeTUzsV9hLw5Xd+hh6j30kH
kGouCpm25osW/uiIX42sP1iBfo/bMoFQUNtps+D4vxdWCNVMoYdYuNnxM/S7c+N0lGSwO09wx/4D
xheeYaz6dTkD1BWmURfzme+A0pvp+t0coEJaLPQ54lRWOr2JAbYyBe+zkY0z4FObAjOQSKFIuRf0
6qSRRDUoQqO8NkzHf8alseQ0N/63icSVHKo4GtQvKXCiy/XoO70GPVOC0dLfX0eMQBql1D49PxkQ
WnaMmufiZ53wZ6+FBITb3C7/0Iv/Uu6AaixMczgC36j8MNoJ9zcEiqqwBhDNF2hNznwZfhNwSlpl
opMNRnXcLrNj/O9j3YhpPyW24yhucPPHcFz9zQG7qdQQO0Jy+HnSyehD9UVUAUzqsU+5ItMPsOFZ
A8KPsIg15XeqY6KaKmMZbEVu5PL8OxStbaxhLjvczKNvb5+RoxDENQYF4qwAOkoV+wepnY5LUy3O
uswO7HbZe9p/D1W9JOnun2trpFO7rrw8Q5uZh9tJuO84c9sDC8kHotLEHWo/XmpIMKR7dKkm3gq4
Kql+ikLBpgJBDnwCY44SRkwefsvDzbFD8W4XiCtDYbDdzfPTMGXQoUh+4/ABICr5zI+8UoLntYXh
oUriq9d88EInQ82h1OSJiByAjXcnYbjmhB4tJBOF5PcgbB5MrSr8O0JVuIMIdvV0aem67OwyUFsz
NB1PsRA/vbbsHX/kWKjCw8yCPpEAlTW+K22HYAj1CPHRUgMnH/8QqMrmRBnI7Y/lsMG4Tdq8T8Di
Tt5fG8WRzvkJS5+TZV/z8Hl0EBc/q2jJk+pppaTcviBIUehbGOi14DV5t237lVXkZ4ko2v+u4/8j
JtUSiTU+l8Qy3/opBzN/kwjkmbQZ4LwvqHd0wOQBCvK3mBMYDc8xp/GXTSlVsacWXK/W4BO3HQQb
bJfjCUAzgfFC7Ecyinme1lOMY4sdGSGCUGKjp+8Mc1B6bL7xu0Aul1UZKMEuvWWADZDbM8w0gjoa
tDv+aA6GS0n7S0IXcE+DM0TnZLVSr2pQaLKiEuIvhA7pTO7J0o5WWmB6uO9oh6Z8zUwrGhQHS8Vp
ek0TJoQ9htk9H/506u/cd86bwk+UzOAtjdZ3PVPNd6+Posl1gBRvIzPESAEJbfPNFamKxXhbcnBD
UOPpYDo8mE1OULD2zDtpB7hmMqwcmYjoxRho2+KULdW67AUwIHPMbvFBa4UD15fgL8x+ueH8E52h
a5MIrKMRLPCICbDsoTCM+aRgmVTxPymyKrla+35vOuR1ZQvr6KqEW2hXlYBXzigCcm4Acbsqb4Sq
Lvx/iEC32kn9BsYsUWoZ4wvug9a86Td5G9xKyWu5r9tX5gUBz0k+Fe6ahXsNQaAofsKydxS6ZkoL
Xcece3FgYIUrbDrFCm52iaSjYKwTSS0R2wYJk6zjvJxwy4OoSQnuUEdfvijBnzi0hYClazkZ149g
yHIUD3GUSJnf3Jub4L8zMOO6OyhyF0BeIfduajC2nUMSSxd20N38ZoDR6p6dolCBCDg65bcqhXIl
bCPOqiqTvLdnybR0vv3TqnoFfHytnSaeKKC91641TdzSS17qy+4wI6wnd/53jUGSpnKh4nzxfyuW
1wf8soe2v6AgFRt484MLyiI2W13j3KHUif2Cu3DlKtBKk83FdvIIpoh4ZCRKpTOLZIvFDhwf6RGE
G1eICFjGRJQ/GiYQgkzmhtII5O0e+KyRnweaqlLz6qnsSLK3ZzXFrJj+GKzyHYvl1ZLLnTC2ujLW
kh00qkmbbHXGzhR4XEk71gFZtjbp5tmM4GWrAbjx0nZfFVAerCzNTaK3KojdkPjE+Kcj9V2V4KbJ
/p/5FGtq0XjKvwOtEuVK2X2HS0L3LFG5zvruHptTgjHJiG50jb2p6R5TtJpeJiAENs8l6+FAT0u5
mULxGf6T9YZ5Ue0WTi6xLMlpF1C9/V9Cvtn842gtoej7BSSzGPo/YJwVEW0Sem0QBflvFJwoTmO/
voanVw+0rsGfFBtF+TjGtrLenjeyNUPeFtyl/nCRrWWF/0cHglc3VkAp+t7BFMalY2dHflW8ynxu
QerAMpqhIkDqgvR/GoT0WZ5e8QnO4fvO6SWyhDI7rExEYwM4b6T0nHcRTQhTh8vqgJrxFeZdTsF/
/fwLkWb7ry7LeBVLmWipuBeHM9DNUlggSk789kA+gi+OzZoqBMRGxzAEf2ym0dJb+EZ9NoRK6QrI
7lJwlwTO+vkABmlhZyt4mPe0yWGVcxrO7Oa/XXgBQv3lv1dASQmpJ/riNO9VldPJ2Wb2TQdskmTT
Z4xfZoLpzYeQKehcW8WnN08Q9fuS7oZJgNc7qcMSd4zXXKHB93fARomMvybYLovCzJU+KNqHFXGj
usYB7HbrOBfgtXsxzFEyOvtuGzeqTuCOXHOl7Hygfn2eZpfP4aSXFI1cjxMz7khi0iiuBwTTVS/R
d3A3+GXhISS7fek8kqoAryth6Vlv8VcYrcTuewscu5dtLi3WPx1KFkLF2r1OJZx69DnwB6iJS2HT
X79ckiAp+2pzRfxLBW3I9K78AzTV9g4NYrJ9LgmK5tizGysfjDVKXtGt9Tu2da5s46KOIBjEDRE4
s9WiVDDEUWnZK5MZllK6G5T123+l3qQylBKTYsZjXnq3JnUkYGm9YOBPhAcb+RkCMyJXMHU9uXmQ
LURa2GfC0pIHNHVus15Aze7+DKRF2xHCBEISDYSoELpQ6HfT2G22qIz94HO+Y/7U5jl6+uUYjt4j
y6y6OxvczdO+/KXESHVv7aEROOxQVS1hU0t3fc4zD0ZMhEqeB77fPk1ZXUyvRlj6KLgzaMqGdx9N
4vKHJ8KoS73FaM1pK2HZCYwx8omUUubX4JTLKCnWaOVnAYiq+LQZti/aB9lF9ktga+tTXq0hRFCx
c3jB49v8Ppqvpm5hHCEBTIDOHOLGHbzugWuXHA24IPTPqzHMfKCtFJ/H2hEwOW8ZZ49GTFmkbo54
pYeCGN3QeIh2+lWjqye88gU0i+6khYHiZzjXjG8SG5rSK/xCgFkTwBb0UncWaWU5cwVCoYtDz59c
kvkLzoUsse/QWwz+iWH+Z+WPxRoI8d7q8w3Q7DMVqqXh/LloUVqxqN3E9g5ivoF2vCnWtRqSgAwv
jym0404AXjThLoo3sro+r04B8r2tOH5ZQpexKoRJuVmAW0uGd8ZHxG6MvW3A+hNL/DleHcHAOUE9
G3zR63TebGCXI5jGAWSAtNOs/+OKg4G4sj9IGF/cPY1zbSNigUysz0yHxYJnQL3gbM+WUqAXzoqi
c+ZRoCBySRZhWlcS0bO+EEkJUWDfSB5mTSD4iq1o2bZXRmQPkCt+XgZ0CMGabvHCUlgxmaPeAeKe
5Mx/Gl7wPEP30MHMEHr9nXJpC8Ukgadxyx/6162UJmi8VkIEO7O+Wz+kV67M8Zp1viQif+1ugKKC
qKaduMhVzAJUkCkT6X1s8EQ0FlabmcFXtStEX6+SsDuTLOzsKGPNMj/j04zwOAPP+mwqF2wiiYSJ
lKjEUtYBMwotiiJBpDUrKI9qX9Aqtvo5in5zbYqcrmSzIHiTqNbQmlZN/CG8X2dnrcbjkmuRGUxA
RKgg9V1YnVAhha5DjYy+02k3UMfl7CF8N69QBuVnVQWxLee8Dg7HFvh7+ylyleOzy49Bc0JDrdrL
J0Qy6Az3gGJKXWzw0QMxIjFQP2mzSUJo2nMgvQOiIAEueL8VIYZf/yKctZs2u51cuJuKEzdm8Y77
mnjZ/4C+EoZGzMKAk7aVJR6oUtFdd7WPKnd0eMyuRIeGSvIpntTU1n+jNZlbIzRlnCnzVKpCBzdl
y3MjqQjzd2AldZNsgS8XLc2/Kegr6WiddtYjLFnbn7pINZxpj1FuPWfYVwCRIqRLctvB2Rbv5JxP
RoocIKFGHiTN1P6ZkLEJuESUjrTXjqyMbV2tYFIZLDC7ITWLNTId4qmv+RVN1DFEaswSjpIl2sSQ
hGJ9LstvWSo+P2HzN5CsXbu8OziGQrn4dFiwwBjFeXlFnK8Nj7IX43s052zmCTuC3Z8Rlp1o/oOu
YDlVTCszJnVR29yD7gHCStFunuRr8T+ZXS/lDmtnyMIgQBSzY2FfPDhtsVnbsh2dC+j5jjRsuTV3
mJZe9mQQk14IhcYHoeaHHAXaXgUwk+9mkyZppxRaL789FMrv9EAuNlnfxWjFjlrIcP2e97Gm68hd
LvflzpO0m4KEeNNYYygmD2r6i/h4HBTENp4uTtrT5m+ICVJ7us5Xdk6vh0ue1+isjexTdvIso+to
2hdVSU1sJt3JZorbhmNoRysCqNQl5XH5EeRgzK8sitmKY+gJPNRm1ORoJEDTRHOvNV8hldJNbZXT
x5FfqxppWYY7bge6uAYjfdeBy7Pa6J1mvGeVR0oZSHbYIiHGDSXFHB8lWEoZ+InPG042Y6+AZaIM
31+yd8BopszEh0gMlKlZ/jjH9vaE6plmPg/kYZq6mh7923pL0HdlzUxKe8Jgtk6005kqyITwpgaH
jEcOqgB4KdVoI03oNUfr/VWthIPDvkMVHsXMZyxWFyfHDzLDKWyz6pQI0p7jaeS/p6KKE1egbm16
WoRSMyDiU26JAItPke1Nr3lkr/Agj54aogwpz4VE8hAGdCA6WpG++TnH7sEgA80i/WsmLBM4uLSW
24kvYnO1J7pU9uHO0/vCGtN1MzrmSGT5A9OlPIHxUaHRjUbpTFHFYnlcJmMEeq+bHpsvu7+xPCPZ
oeQ3ZMQELaLp5F0zzWE7O+LIYijcPip6X7xCsDa++5J7QShfnJnB8xTtSAg7KWBoB1dgRnKGGt7r
ah8B2f2zO9PSj7DH2moXCvJWDwadCulLKskbOABV0XXEL59BJvsKqn0aP4hJQADfGvTurfCNDaxx
0nxLm4Ienb6Ovjp8nM/0gwCa79imSeAfZXGWH4YSiqlx5yfr8LQ54h5hk8IHqX+LZcLbY1i9n68y
N4k6M+pGHeLcC91+HWe7UNy5BGt/mBtnb8OqJrqfGmBMnQWhpc2oAEN656BtBvc7BOFw0W03ZVyi
X+EH3KrMz0l6kZGGv0EcJsOZLnafYIs4cMXWyRGmoS1MG/4sm1tCLHl2PPei8Irjn0auYCedf0Zp
AWtodGuFpaPhx1kywYKrlFm2279LAoHKN8Ss34YD5vqcjO2AqZ9qBgU9RI9QS9m3oHqFsKULenlH
rOqjvM+ePEcSkS4buU4fgxHtloVOOXNFM0dzCSz8SE2H4GxDsgcaPSKMejA1zu0uWz1d2hAekWkC
gMJ2f8WEipy7YxIBUgAtq8NQq97Xz3b24myLFr69ZzSM/4GCbZ+8Y/WKpmViiezBul41Xju1h7IA
9Gn5793fffNsASD9RXshs5ugTdojbHd6UrhpxkMBrEYK8ZI8yEA6SmbiV5HbLQsL0jFpSdnB5+ri
i/mHRHwDOnK/5MKZ5s5VLveLiGg9DF8jhpTwH7KMdlknCr2wwU4rc9L0Mm6khw14MPqGJeLcSj/2
hXYcp76h3fc8Gu9pOfIRrlrMYVuDdkrQS/xQq1SFG395UVOpAV4zix+bhIl9h3pm8w1J6MbBIM7F
srvbL6sCQGdW8Ex1TYpyoSRqvLAqlLfk0NIQ38Eyd8vS7hKx0XOb8UW1tTayYNQhhVBxQgCcMkxH
s2hXEqqb669l7NBV5xEVg0t5/HehEt+ER43/UuX/F6q6TmeMoHgKyKG6kFhpc+RzV+In9ZLTG+80
WQV7Pb2ldjr3RcNNfy8nXLa8LYCWX9nC1TCy5v2IRWo0CE4VBXw+D+OjCI5UfjcobTMyT8VqgNpG
V8+cEKMTCOjxwwWn6nC5AUJc8GpIHfBOS3QnS10vYLXcTNIG6EaS8kmGjcv57CE9Kfu9Kg0aLkvH
J1MtuEc3CkR4eFCXlBX3iczDqXXQLD76Pba2Vzgexe3JXkw4LYS33DO7GEU8d1VYzSJ/kGO16HF2
41dmo4uIHypE63TSoDqqXNk3mcWUomHVheJtXa/3wEhObUQ2v7snlCJ8Ld194TfiIqEBruyIasUn
qqFVlMtY2EMyccWmcqUv/aXfNXtaNnCvMQudZ8w8JYstg2xJcSn2zZia1z83ZxmsM3wpB+oyBfBA
jGa2jlQw7m5rgiRQ8ezwVl3m8mxDoZPYakrxD2oHe4SIxuJATSMc0mIwlnM+acsXh/U7wbQEq748
KJ1vXNjfOYVjndZbRQ4lzPhQMC+G8bYIGjECkN4RRmftEr2mDCuAvtpL+aE/zw496jB/Yu0HV1jZ
K/lIW2SKXDyps39eVNhfIxaudtYoAR0JI7Hn6JYMkDEg++Fur0/7CKv4To4FW+PkAxUMaWFUZSv7
Y1ciCPclpSXtetfGoxKGp0h2XOtzuT6tmbqZKhxIFDq0bEQpBL+Q+4Dtvt3a7kUzWLMP1VTUDBqp
Bf3PsGIxp8YyB7tFqxny2qmejW+hEawY0L9kbMBid2IHlHO6bxZaEd+kshYpZVCOFTGLmll6BJa+
6Frn/Mpv5qc0dHVImjnhciUpZP4vOi6Xj0A4SKMlOfKnfuMolRG9riiHTxiVHiAMXq7bG36tr9ae
CzWMgEMwXVYPdceKRSvG00KWAzEK+3GF1zAD8FiU0yBRVTGcQzD9nc31TmovLaN3yVckfHdtkQfy
zTGc5f+dKd/Sg34LbrI/ofJXvhzq8AuLcCDEHnVSl0vWPKnoLvHEpbtEo064E9cL5fssP66hKTIv
Ty71uOIQy6HlejDXKYvvIYbpzJ551YW1joxVuaIFMuQzTQEQEyYPA6iHv1kw7auHKmPCIMFhiTyc
pAGw5SYBqLBOipTLzRC5QCsJuOU5aqymO1xZrNpFiBS+LaiDdzzIvadxwGU+J7nDuUTkW2ZTFx/B
Rx4Wu5cLtKm20na1DJLQS+otk4VB87+J6+fc1797gicfl/AyJZlyuDJaPMjX8mXDTY5GGcufc0Qq
4p+Oxxb3jLFj8cGGkgGmJuG8xwh2vDDcee+Vq+1z3OLbq/TsSgyDCFfUrLeCNjNyqydyG7S2WIBJ
qi9DXXzEQ0cw6Yh7x3mZUG0Nj9L0Y/brcC4zEZlMOVaoSU20Qt0AsGGckCquYpcPI/52T8oQEq9K
bmUp47NmWGETpmRkOlBKJQYoCFbKJa+Lk+D9oeSVKsh6FmbxM6ZHx87jSz/4jssN8r9GJw5iiY5r
b5m0Y06H1fenpk8Kt/+EkddsILtDaLGD3nw3rm6GizI/7omRiNSYG4D/2eNDPkLzql5gKACk9SHK
frmFyXmR67Hs99Z59gy3WKwWLeAaNqqPBhTi7ofHaybyQlGSl1WAkhtQJrWo4eXPNF1http1i5PZ
cjtDg3clUDMBDqhVW9CShT8rJv+NHj126vuUxznMBkd0ZaF507QFZk2HhTDi1ANo6KagS1XRLU7c
6Puz6WQp78CLTzK6vkKMlVZMgHWeMGg5dSH5tL4fUqbIF91nVhsGLSbpQmXnyB37CTpe86whDxnF
YD77rqHfHtOUyqp32ibNopV0mwbHiVKUCCABQBGGBrHUU+2LcmLfL0yGiLz+e2uSbwdYs+LUWr4B
7dKUxyfkE8KR0Ygjgre3GFxIjLHg2AP11irTKtSur/5TJxAhmdc+1NGwCgwsrfF5axeLV5xTnm/9
77wM3xyXC2r+95EBq+1XMf/g+DmeGKHTPxhfmvlstt6NlFpbHJSvwX0mrBOPIdmFF6XnJ/hSKgs3
nZ1KLxIs+9x00Tlq7OSKBHRzNC0o6i8FlwSL7Xc1Gzc2OVqX+jycZBziN3/lVILvOlY+p5Cx0yAj
xtdKGLgyh9EnEjoN6z/ysNDWOn0ZiFJ2QpCqjrtIDK6LEBEnNOjICvXiA33uqG9u3HA4seS8VB8z
ACc5ISEgnyU/AXwRTkDJIMS2nunAIso/8zr0Wk66Q1fxeEFB7nh9PF8Cj0wH7PSOB3daqZdoE/rZ
QYzIOXbR/FrRB7751NfX5y+PxxGlg1iCjuTLOXXpl4kLL5KF9eHbJZegX2lgW665hzDYi0S/3P1+
8SH0UiCU7D/K3zdYY+pimS8qIdlqdELPJMdENPWTQ/bjsaBoIy2KDTN+PQzWs/OUpkcVPHewYIdR
S00f9PXb785sMFaxE8giUrEax5oCQ3IWEhF4WnZDtt3rTb5sY5jkHbrQHGunwzwH3AuwJJBRhYje
5ogNtniL9fS2VwCFok+FfsGhVuZR9g7KVpMMExooD5Ue42fau3hJy81Dpd5ycR+O0egv+laTVuVQ
6dwy8goFvOrSuvlgeF/0c6pRKUloqugaO9aE6lItgnAYyZK46t32JaVYdzKfLPcm4bDCDeKw/1+A
Do+sVbrBE+JOh05r8ah8rZqgRwr4MUp2vwnXDjnD+vNBMo0zVB0W+eCObqPIdfel4hkCGGygpIQI
9tgvEZy9KDXvkK3MlWAMZS2XmWd4X3QINUtlgQoPsE2cMMiTW0qWPBQ93IpT26THLFoZEhQA7j3g
sHvQy0Eb5mOyJVFo7hJNmHz8UZxgWdHOoPeBqdwUbnQs1nmoU8tBKHQJ9MZqBKQfzqxGxRrtkCxx
TCeDMe9KV9yiObCiIdR9XqweJ5w3pPMszXIbwrfhRLgZF4tMVZFQaqs/wRXYoRejVvbwjIXP+lCb
stZNqXu28qvY1C0iWpmeSU4flF/LmKsqBkAR+B3l9V7ZjpeN63kMnbxesKULJ7IsiOpwnnqZw7cZ
/tjDCtIcJA172wJoFMq2lQ0BIwmxdF12/iApWRRofVsskFBjEN4kMnxHXPv055pv9wvxuPjeA2Mt
43b0eYcyFKZeWuq0qT9MvvNIrKAOtKZDVwp5p0kbWRFkGsmf9GVORpU+qJHX3Oq0XXv2JzRSbWyp
jOQYNjLtCc7drMyTZRb5/GN+8x4+VpBal82a1IrZaREMp+pXNd8L9pkhAHVN9Ebvf2M5UzWTuAO4
Wn4XfNBLTspscIwG8dn4pNHLiSJZGRXv4WI4LbmhZhneRRLzz90wXPLDV86S0mee01Y1mfz+1f5u
OiSFRXSgJ010izwOZz7VtkKtFXhjs8MsUNymLJzEIl6YPeIBE5UpgyExw5jkfxLWEqCieR06gkwO
k5cMrEzrWX7owo1+TrhSahqaXwReoP0nVEdVQUzYrHnXSGOwPEhm1GN+9vVuP0p8VgWJcuOYvDLi
HE0lN71INJqZ5kBmolgJxWSlBm+ucDypZ0mJmQymvzBYOrifuMxYm1c60gq/vhmQ1Bb/Qo9ToJd6
V0x1+Z3ca3esz9p6loCO0GMGx3+qYT3WqzJcjUHBdrvKbtkh0cSorROEvPTUwqbaqeHdSilQKhj/
pOfYmcAbNkakFDeBh9H5C5MKM1FJZ3lEuKkbyyBTrrnStl9z4/k9QdxPtLbZcVUjG6JYehDMwBxi
Pj+eci3dZJN9yYQI44c9qJQZOvfWennmZe4bF39vksY/WUn7T+NlPjk2AjppImYD+GNHz+8MJ3mD
Ch183FEfqBNapoOZY9C41Km6DArTX+XFIVqJ/5+6eZ7oqS9E4Uh4B4NoaCJ6NS9JqpOMveQQICsB
TVTdgymp0hsLW0/d9W16LmcCD3bF1LG7fW+NL7dn994nP5/GaXlJluv5QEAuOU2hygbMiLXE6tYj
CmtKYFt1BrgTkthD+q7PSC0yq4MDbSp6k3Oy5ROTYbNszwFvqQXZgXhEJQ9DEAgJN74FX6Jhf9iu
eJgbaftToJOTkAzFb0vsr6e76R2TWipnkV5KEEpReP8LEzQH7Ew4n4teB+NSQJ0r0IF469QaRXdj
G508UCU6JgrvQ7ZCbfkyEm2L19tf+S63Cyi2RcY8wxbNc2nnbvV5LpUn44ml/oKv8/fdu79uUu2u
53a/tm1bviQCcF/odQYEvt0qRE1ffZgsIYP0qv31hE2g088pGEV4/OvmhwsxBg5c+tT+NDc+iLl1
PmMYfARHkOlckGoUMzH0uKCz3q3Xv8QzpdctHSPxx68PKV+vKNRpKIUlwUt0yH+trjl3lPHWUupf
F/2arCrowP0zDmRY3GUzcd6YRsdMZ55F2uwagvuTyYJ1i/KCq3wXfCPjRDfL9kMaGDuaVmU0mO+w
sDyQxAeVjVc9vKoBYWoWcrN/DAp3bsUekiEvjGLM/CgMnIxVNcX3SNauCBBBCsrcqVs1opEXbAw3
/fclTaxP1B5i4Sbtq7STcBLXGQ2rcju6CBrPs/LTi+KpQALLwAyXfbZTBf1tDKTMfGgZSkl0Rd1Q
jjRVTKntzWt88T6mFocatp9Uwh01Ddn+I5y2D303cXLF+PCeVTvTSDhWacBMZQW+npH7S7ZDUCCP
MBpXRxuUi8ecTxfypG2ocTBFaY5phtqaj0zEehSvv0FcapIIP1esqTpofsknP6vR+FZ6b38N050R
Q9FBscUzCzgBUPK0nX5/57Q44xdmlUDnoVbMLheIRz6ae0vSeQqIUAo8lYxOrQn7NhsLj+vIAFA/
MkoMeWBTfr3Pybl57udHfxXQKfU7g/0oFiwHsF4d0wsvmniayBZaBwJOEa30CK/DAJ2knG+KUZg8
p91iOnrFErgUnd8sUBR7j6tISw1KOmZ1tRN5q5XiKiQnu3onJL1OvKdG3cm6EULvFbSPWLxuWutM
vpMCaD5VrB528lburVHYJT+6iH8ekswYQZAquSoUX7TII87tzZjp/amnbFbuiMAZStxt9SmWghts
aYDVIwExZXdNytR0H2iIuWFeVB0L3GK0O2KKosuhCm2lyXlWBFRqHmGBhkNhjq4ptAr6/Ro95ySq
I5YmfodVWm+f0UrEalU7klU3Hr0FN7ApPR5d669//sYLeVr5X3cUd6cV50dso7ipyW9FMS5+nnIP
SB4U99TS+Txl7/hKdmMe41/NRSaHAhL84cW/JOvHamfDBx95tqSA2R6JjoRyedQetlW+JwgzZ6g1
DiACqE28kK1pNxSEoy0LU8e8gv692Q96lL45gJcojqaAQrcBhQi+mIupcSRGivvzmuniSCAqHLcn
xDgaEz2Ak3yt44fScfRXi2JUPOR0rDxKWjjntxpITmWY0PgQ8HmeTzi5sfsdTKzukNmrUrNjsnu3
MN2txdEPFBfbspqZQHw9YFJwedFpYvQoQM6q9gF41v+3sMV2fxE1VEQt0/+igH+Mj4NvlBwqOAjX
7/XI9ghGgz9Gt+vm//GnM5jOXyNUe+MDP79wu5AZxSSAxZGzm5mb2T4TlNqn9dTDKjfmyU3xIlon
JqQ9LdsU24r75H77ArLVrbJ51Szp0s2f9+ICKYE58bC3ctV7HvreS6MwOn2xHK/SQ9R3NXx6Stms
OEax6/8Xn4TYKHCKO+KHqJIoVJnomDwtGxcLQIVYUOF/rXl9amHK5RrhMkeQORwZ9FjlTVblZHXb
iunmJpCsBRBkof5e+a0xWQw7hVA/T9KuL5EMVctCizrTN6oZuyWRhbkUdlO1Ty7qpt98+1rx16lk
3bVdrLURGvhf+l55jynq+x6luhA0P7PoftgJSkrnYpc9075+kQnGA+eUgSRMjxQKv/vHBq38nOEg
8ua7iibv0jGxVgW38347jBcAnnMtyZRwbJuoUSKMi1nYnDP0BY/vOv/DkYTESjJxPlBfkia4xFJ5
AuBFfnliCJcwGyeS5pvYjfsAvTbUTbavk9yqc1AkF9lpubTCdsQmb8IsLBBdJMs1N6ssDTDbAGRF
jrSGyD2Zb53hMBQg+67IUo0Zs+7e/RNavdQyNNX4NPu08rLYhutJXZiPvSGsyIz0fU5x4PKAejRT
CoSM5Rg4lh4clTQs3bZSBUBHQFzmKBxvlMq9CBfcjN/JoBjfVW7cpjFFoJA/2onUW0ZnKtXQ2H+N
q0U+iGJjj7qiurzY6wqb43ao35BaPVhTrwr+fXQKe1Fix3VEEp3ELVCGobYK9mfMobO9Hf3HXcWX
MjKI6q0DnVj50laBmWYFkQMNy3plWLI5/UzLVlL53MGLOS9B3cAfiw5LrLn6zcp9dM5/2Sheoxrx
RZw6e+qAeJdMepccKydEzhrw0m6ngS9Y1gWNkwtdO3iGPC3rZtnhSz46GY5QXID/fvbdO5qPwLCG
BQhNxv8dNwlnq8VO/HQ7eVjVjH8y/4Lrp6qF/B67CdTKskPAlhEBj3O48pvrPriD9kzSrvMzP4EK
2LbSOJhBKpBLi23BsuBcCzPI3tWrPeCsuAvF71XukUe/EKn4W941ijOU4LkWu+ITg6N1rFbZnC1t
AS2pB0vuqLTHpwwy5uywfA4vboWrAPQmfZryiBpKMc2hGe894BkrxGyHhNDvV3NQ5stcvkL+/Ct/
l6Jm0wEjZHo59MOCg0sSwz+/iHSIHnTIOpCagi8NQYF9EGIIIPZySNhBQ+zdybpG0hemkMXcShzX
MQJVO5sQqCYxfyGJpyB9wU47CY6ICPBf/YT4MepLmNA4hqSZLACenq2mFSMVCD+sXkXsj/6ZG8/t
WLmT1ygseCka+0kBwvY+GZgppsYb/ezDWC+/ZvmNgikUitJzhL1J5qe/BuzUvt26vSG/hHegoeiu
A23Gmhp1RC02NsaZ0HoEZd8grn7xDLQvLmv5m2uXY+N2majxszWaxLVMHd2b1X3iFeehdQSb2lan
EJDlIHb5D0+ek0IRkVoSMuBgCKzdIPi9vZNs9l8uCwOkKAe+0GlDiLvHD3sMc7PitqS39r/s7lti
y4AamkjcFX9+PEaKxuLHeB6Hedm7/U/byVTWAT6gaYDVvUyTfkIrKw0mustJAoqI4PD0DVpMmXh0
tSqw/p3NxhH859r9AcUKJXHiIs6oVGN4rmEW3o/QPhRnTI0XcFP57jO8QVHsMHYpbr7FvOb+E55w
Rk6efTE//YIYa4fqkPFV5UogH5JSQsJ5fTUIKJV3xfH6Q/MZiV/ex2PjBwg0WghefAja3HlgYTiE
+KoZ5maYkQRodVUeEyIT2i7N4V9UJtUnLeW29Fscb3oxgjRnCEEh6fwoRRO9+CH3cbVXA9bv5rZZ
rryS56J/hQAyvfJQ/4rCJ6emVdDBrQJ9BrRn9cRfYH6jlunmDOO6lYdd6IWiWfdSbhC0NFBL63ET
j+nYM50SEwn+SuGyjLokP1IfuINFGcpJatkpbfWbnxLzNTZFKgnmJ6hxg+sSIrqiNx11I6kefsvm
pfdWDNmX36iGQnJh8ipZDHtm+9fJTMtk/Pd6qV9WsetFeX4wm99jB+WSuW9i5TKn52gNdsP2NeA9
uuK4CV5XgJjr93rjlu3WIN0O1GQklFhAsZ45oreXd9FpIGq2gFIDyylFYB8fAPLcfcVfoNkfOg2C
esD59Y9x58++AiAC+OPhAh1S2ApvMNAaOfmak5OOD7Q46LVISIio8eQvFKHcRwM/CbGC1sLVsnS6
fYlUdNLEMTgnMxqyh6znnhPbLqBqv1zO22x9fpP2da2B2nTxbAtRg4Ur02KtkqI0lxGOr4gkWUuK
UloI1we7/PA/4wb+DWBOS/yz7rEEBagzF3FwFE3OuMu5jzR+iYvQkeIGpt/zeULJhkZQiB7rCwT0
KgonMGviwLmvmhyzXEyRJMqyxxPX1GYroPNkpJajirq5XDkv/vv3KfI1vJFmBZ+/CZjBemzo8CV1
EBqLDOlwynOb6vcrtta5PrGpre+mCcsravxKfp4GWWtPFgz4IghuvrM/TmAKTPyLTZczXuVn45kp
3CQ5WiX+TUwpqlsZoJt5yWpQALl3nLXbGgE26gMCGIIBvtavBGJUV3zET4ONXbuf9S5+P028JhxO
xnu9wcB353locvrkX/VJe2rL4JD9xizYEd76qhMMdwyhbWnBX1jal8dGwuIrSOYBTdB1TX9SgzNh
rU36bl3OSYHFqSO64bD2K02Rj+An0NSBTCF/tJONwa6fqFaa+0NL+Fg6yOrNPXxQK/PRnl2XM+b5
15wmJ0IqsC3cfuC74r2/Fui21y/m7NX3RsXJni2uPixF5xV2DAETlHo71cZ9dgtZNfMCIT6AqPeV
jeAmt+ysGw2GYoD+FkNehUoG3sgz5gkbbMzm/Q6yNKGeXep6gjVTamLY7havD5f0Eu2Jpp3V+LOI
sm2eyGHnEzjiCwWfy4IhjRBcPbeYzshyQdU+lhEiOZikahLOdW66Nn5EtXJqfQiH71ez2ccbaOsV
VhsJTbeVcEk15K7arOTIOR4wMZJgnix/rctB/vz8/B39hFgCgKGSFwI2xkfPRFIKWrU9+vFaXuNI
Dn6uH1kgzsF+SSOsSNYw1p1vv8SUqifntSoc6csLCVmHElyyhoelGrYWhixr2J+iDhe3oQoWn+KF
r/iaobwkwWF+uDPW8xh8ZgePeFtoGgGuLoCo3nokiNJ+D8TyHIU8AvEeg/JbBb/qcSXH0NEEYAcC
Sm6S+SAg52O8rjav95Tr+HNGukCeN3z3UzW4QhZW/rMJmcr3N32E8sYdBRoxGjfM31+rvTAIs8qr
dptoizFcPoxAnnh3eIezy1vmqDsBVCitGfyxdrtXpVYiokXw6qiRd58MZ1DYS7jovtu9ijMWaNTi
RoyLSEVk6Kr7ktZnmzPkC0I15he24H9uIp4liyEnMzcjOWRZOY2JWESPilHKVf+1uABv9HuucsLi
OABl9EO/kfTgINsVOQi5ykHmE5B1bK7EtUSY/U1r22bOQx0vUvPEtM8XSMPg/n7ujYbIlC+Aqmh3
xcvOEWGWLnAdLLB3wqZ2BGJ6JTT1gI//x4IJmM1VvumnUVFdvBnGUbxW9e8NYHbueNDDzwvnJecG
q2RE2bXxZ+as573pGABzcejGkFP7ON6W2rJ1ztMiuvYhpizSYDotmSdN/UniuJtxmdYEiLfohCwh
9Kcj+6nad4iRJF8oaZfUyqGafR3fLBEXbZHBw6dNzGLlVc8P4YAnhNlGW5k7960SyBMY4B9/BlJg
St5121/RnWUP94rngaonIzo9pjPK8t11zZyJxSrNjmYzfFToLh8Yx2QTAm+eSNWaW0by9VRqO6Rp
93JZK7cMtLzolx9r0L+QDKdkgqov9+f++Mwbl7mraCDyne1dEnZOVDLaW7uzQAbbEXPRtLOsKuZZ
a9emEhdtDR6nbJRDroHDyqh7/PSq0FUrPlUHSKFjK02HmeZTAdOE+HWS7pAKcxfVj1bvOyuF+FS4
kit1y6KAun4nG/Hm9S1hULsVBUvVNFkBxJNaEqjLaa1an81hTXESg0Ng0mCwHTqtWTIDcEj5Be1f
lwhqprFQyWEAwJzoxmycCnUuWgsUK8+pCu7RaJicu9q/ijqU8YKGRz7OPd5IQXf+Z61OUfP5Ubce
KKNGxAg64N7OJ7Rtgec8672ZnJ2iTBKNww+7mq8YMr3EEfyexRYtgbQEHvHdQ6XVXhuHxqY8oqxm
yrLIa0cXatuoTc9IKPwu2qHxYGJTox7HcD+kqYiOxj1FesvdN3OyniD4sRAYxO8RONavFX2CoxtV
zpGF/2MHHLTnSyNjAeEFXSYjkJKVPqcyLFS3KRPgtmXDdGQdkH9j1c/h3gyEkeuxqRMDtvbp5vRZ
Y5oBdEB7MAYORPBRvpF8qtPVuZrDJ87IbYu15hSFvWWSYQ05qUfYnEMbWsYDrJ5hkIHsclCvLYxP
eoI8Tt+hkNfcKGwIKHWqxd3+DXrYtNqGZgXed1Sph3C14+mXCyhsXeCyjOs0k6E082WaRPf9c5Vu
2ENfquc1brqfQzUpIVC0zkC8ndU0S3pmbQX3gUSvVLBJ96Nt+Gx4HPpRhsu4AwsmqgiiV1kz4aDo
dWl2ji3sbPB+jaGjO1jQ22mlYdh5s4/S9aLbVabb9MlcORnLTIIHmPa2Im1ZzSWlA3qvjZbVJOYi
CGTQP7kY9a4+Wg7zkD7KOlEeQVJYgvm6eT2crbSiWOzu7usPEJdahsqP/KSHlwVWA2X9RNCXDTr6
LB9J1wdD2tHBqXyk7gKcrSer3eCWqSeFp8EPlbhFmZ7GcXTJPx1sPj663ww64OmWayCvKMhNxf+3
utdwIrrZjtC65Y3C++RU2OOXt3ODkR8sQl5q5HAWbgLUxi2ojRPM2bMp+1UfCQ1FrmOKNsJ3RMO1
snFns1xOWRCmK487vYcGzcqOF2BXUIyeaVaJwP5Pa46j8FH0nYGw5vG5U3c3ZOql0BxnWX/ZoJyV
re7HnpCE91muFioTG/q6semhC5yGvK8MgQvcvn5Tqtmrcd0+vWXnn+fudXvfWCHyTcs2AeyBa512
KXHLMrDdTGorZtId9OK3sCyQPfbYpLyRxbeZIay66cjY42tv+MDrAaaOPgGK4mnbaLOmTEQKWiPX
/LktbUafmBld38PZMwtiAvTqHLvV8Lb0UmzMH+NeAsyJcw/QfMhuRe5qLhRLzycFeqEOhCS2/9Zw
lhJr+LydofN6l7DA/bJxxRNu5npfQtmC7DFOjMh65oGZnhH9i+v77M2CptE027BDrEgaf4QttCV9
zlVrwJs22WeqLRlsohQjOkxiuAjy1JefuJT0sXHWm7Bkv8U43blJYPs6wJtJmeHftxxmWr/Ouj2G
QylRzUc39cposhsI/N2MYq+YNY7JH9PCM35+iGzIHinUZhazqFgR+m7OfWRg8h2HVTQHhTTenMha
Ph7FexIdR08S66foUCYgziCu6l3d0q4go33LU0Vpd8gZQHG4yXvJxhm0JZV8PcpJO1TEdN99JMZ2
mvNXs8r/9Bvi3GP2aZrx5cPxklEBU+YgCXtfurpKjwIr2jrycXcMnU1vrYj8t8KFWYHQA8qnTvjg
6QWJuxmjs0lWWiexwm93JGtIHQXf7VzT4wk83SNJfHAM+FaqktJ5rKbeOhLtPcVSY01O39ADagTt
8vmnPOYF/DEw9awAJBWLbJL2AIP2cH4cYh4qpanfrhE1+JzKCgqs2nzrqGJQK9M+PzJONamnALXO
Oz2gzS6z7w0hr+5q7S246restBGA2jpxv9M6A2RJ+3PK7i86wDlz68ObVuVtQnwAfbtoEtra8YAE
g3rYgMiwkvYNnjWn0gyV2VG/bSnBLueSh1LP3V0Kf5uOIl0hCVyGXqR9n9dBipY/CfiATbwEn/IK
GFH13TqjypmPQa/YI8O+l7DgrZHsDuz7l/xFTuzJh2HHenrDSp1TgmbE0tYLsjhAfRFisH9pJb9T
X9NqPGx12duYTfCCNHPdWCJ5sf/LRMC5/kQfoNeW29/0GA54LK7H3izZYN+RNkwig7FNZeF6EO1J
HoFZW7xYMQJt7YTL3gRelCOOrUbI7DZPOswjp+vRSPjLub5/xJDO8mG9DvAOdaW1Ccuv79pf3txb
WC0vnj2xZqNWHjnILJfxZP58DYmZUTvFfEMTIyumUd1ZHWuCr7K9KKeks0y36QDhrBSHDDIwaxV8
eIus2eHsPa7RgcpplOeAtcInVNQfaWL15xaRV03KtXhP23RUDKKNQcemCsO+NHzP7Kr8X3grQtcm
n2ZfnEtbMkTR4L9VF0Sd53jKppDS7Hwk6ifDtKF4dSWuGsuZOf9mfFqsB8CGbaC93YEMT5Dj61gu
lgJR/HtxifhGHas8DOfi4dhhLLcB3lbBHTZhFOjw+OAfO1sH6X//XuaGZYOOE+5tjAbT9rrXUXaV
CRiiiNESAGTUveIqPe6O6SCmWRUtsnp26Qym0rzPsOPUFYcoBhRoO+82sbtq+Bc+kuBof7AjWo4o
2gGVeAcmSshapB1GL3zk7JYZ7PDXLoXwzo+Vl9SYSGc4vgpabB8t8nup3glFSiPT/NwIEzl7WNtM
8fHWIor8GDHmrhYUGFEv996sP2KhqOZ/vkMvRvbvzqOS6BQ/MSAcZ86m6JKvN0XnI/cSlBBEvqxX
rcLW12/CWRtQHJK6DVKNb9K8J3UJXTjNc8pz5ObAdBFCTgtRAyMD4wXdsWl+Mv2niaViZgJJZquj
nB6FDwCT7XakaHNBfupaIRUSPSqfz2qcipImwozk6sDE9j8ITUsePZgzrUFiDJGW4apr1xLNf7+h
pmKvipD00DkpdCwqKvz75wq2N/FtOOUEK/bG4gnLmJAJyf0ITnzHB2Y57O/0x188fkpz4k5d/+SJ
C+Xu8MQ6gTbJyJMiWIAuNTXrLc2w0u437+rXBZBWzxhmPGQmqcNwkPefoasumWbe96/XEBD4OSKs
AjwLDtIvBDW6Kh7wdFlvRwmmh5BJ6K+MetmlxWmUkeJIcVyyykrGc7Az6uv5imNdI2uGuttjLclR
roK17n2sIFI7AoJaR3zrgKuSHV20fi1LHkXcgnQLSynsvXVh7Xobl8lrUWJhHoOli6o33lVgFUjM
hYFL0ajJmyfKV+LwBSOYeUNAeG2TX7BCETMPYJLN0gF8BiJ5vi6labE0UfHgJGHAG+SZ6kpmdved
8g5qnWVWWQMZ21IbY5EXviPPNhDjsfM6RAWdqH+40Hd8EEcNrYOZONAiP/0OwS81ioGckGh1Dzl9
shNqm51lQI4m41+lSRCp6ejV7UR45WWgNwbCC9rp9xUrLtGgUEqqjwZkY9keHQzSv+wMR2tXXbs7
zlaKg51Xj8ZNQzi+UzqS/H9fq9NPCDQWcU//TH7w5nQw9/h1TmYHTdkd7OrQVGJgjXyxzL1D/POp
7Vn4xuGt55DJFvicT9dvxA6pFfdEWx/B5CBWiJMtF89MFc+WpY4KDpCvvY2WeQ0UwUANT/ZXBIZ1
Dch1qPZlQABmzVTYhKrLH3kq8lTxVh0BZ4eAh8kdnQQZRqXJhWnQ9moLPbmkwKPfhQa9PtDjmoGC
opHDM69CjzJZKoc0DBg+WpUDf+kJLZyAIn6OyfO1jzNoAnDwwDWWC+08fsCVPLnygsG/l7Pbbs/E
ZBGcSfz1mmZQNB2moqNCMqzyVkSCFefoa+qPi1smLN0i13IZBJxAnDaT79OI/fNwspTHxTeQ+19N
Ip8fNXxSkiZ/AI5fKZvO1bZS6C0+rL57i/YJfHKxMUqU3nuiLQ3yGYwDsPkziCLZ1Cxt/oHOHZHS
Bv2Aj/4ETjfZNtuFcAFrwiEHpUBf0a81cU8WRnHu6gTSZz71kIaBM+COCR3+Lp8r1zQefWNz02Js
RFENFyP906CarpshknLUyMYrcETd2LprhulCDaazLqvrwnT+hOUzR+u9zpz5JGRv5NK0PvF+UuK3
okvS+BgB0yhifmSEafvpjha/jR5RpCrpoi80A/8YPKb7FE0QSbu4zo6Gv5sMZisAGd08/lwLFGJG
2wN/j+dkq/3OgBWOXi+Twn1Uc8gcbW8MlxUmjp9S3IlzqXI5G6/FJtfPIhEBYcSdyV5HhbJQQ5Hx
J+2M+KXqiGmopQ++uBlzViPZz2ZvpaOv89+adc8gPUzfqe5bb8JlQrN4QcvngcFnLZPhTH0Cvv0e
XaXSdbOfMWLNYSX83FyS/Uinu1PbdFilBmJNHwDjogg4cHNaAdBSKkAG7W9/pVHP8JVnPZTFcVzs
AI5czYAXxzA4LoS9LtFbA9N/OJ7KRYlQe0wsyNrFQz+bYbfJuuXC9SZVQlWDfL0I5E7SBqI03v6S
80vKIUQvOsZz5XNWnVYqZQM2R23n/U4XOBwjqVg9iQcyOnq6PJRNhc9XIQvVygjCh2JA2B1OCvaP
GPW1/pYbMg8hw9pE8UgWspJN+a/SpYRv4cVFGR0Rcl3lnBzxopqtyQzDQO7b9PFk4Kd2L1Ln1iFl
qvDZQn2gk8jYJLC5uBKWW4T338fszuyeWAiLops0EIaa21UkmQ+f7uoT4iqi3aFJp/nfNiFhI9BS
Lxm6qOxCsBLJLRM4Pg4l8iBi3djX6W4seG4QrOeT+/q3ozpZi6XmQL7Uf+MtuLncZFRlQ6hKcZYk
0Y71DpXmuIDUFnJfsxTR6/IY+aLSGvZXVMv1f0s7QHGmCtRx55f8a1lwGfL7zJxbuDjbz4vdG81M
r9K03BiafzHvn33msIKbdjPLv/XWZaimUWy8R5tGyys49TjZ3PpOXxexJ0FGisid5CYTSMtoCoDm
gqJM2+WT2oy1Dz/ul0CqF9pH7u58rCMpAv68IvCLBM6i4acufJ9pG1hbu4zBBMz9YhujuOjA+3Ew
nGMO8QIIePonjaSAWNr/C22UVfMWy6OCaxYtdwjmrn0vMv6u5xnxshfAl2imyuzaWIjkqiOzUQlN
iqFLHbHgP1QqfaW4oXN9KEN+Q83aDS3yxtweN0J5mX13au8SIA88R+i0nje9mFAE27kTvycIlXv7
ojMjF7Ssz/Iv0e9W+BGM7qJka7Qrwws/X0hJwgSCspI+ds0dyJPYqul5QUWBPwjvOR5DDzp5hOlV
uXRZzyem6OTx4H7S7lt7Cro9K2+ewsf2ucl111BRPY+TIPbbSfIzih6/DpGsqYQYA9EGyLEjAS1b
PphC5pY9QxIU3e3zIxzI7jlkBbXE0kAHG+/I4uUscVlM0g9omzvzGF5jL8A+pTP1FW7i2wsc7qz8
wM/zXGT2HOGSH5yUMeQAUhwq/yKQP9U4r/fNLg6l+S1rqwTwqUy2CVWpQEPIP4ck7rVFXnUf/v22
A0y8SS96PdVy5fw+/sYRzgBsUjGhY59PBdQWcQSYfuVA8HoKt+2eBrDB5VcLB657LHA8ZeeAg3fH
EcniK8GVwuX9/veYU183D/kIW7HdZ1js6LYOydpuJUXYl+k0Tw4HlcOLH3DrEjFGt6kRDDm82LDN
zqbN29wt1iiWiISCTt0agBPcTtbrLOo2/dzPCHgGkjs+R6xssNLHgJtLZG+DxmN557STVxKXPev5
U1cWKQqjQ2cefFVOOU67RR/bUvWGWVgCyoWNN7QWT8/scmejCbaUCKp9HXitzBgkuKNxIYUFQkdi
nVY1cfirrmuopxfzmx8skAhxRm6bV1aLZiSA4UriJTXT/svR5x3Rlm9sqecrBGWpjjmVHwyOztl2
dQo9vzlvXLPi8G8LXqOKgaumqgRizlmnW4At2LWtcJz5RmVAKtk7eNwBDrvGfk+hCaoWPPqITiD6
sSaRexcdNU5lgKh6CCQJkJvOUkuznXy/HrCH+GHthGd9UDVtMh3pTyCkXKUvq1cCQdJWtj13+6QY
L0Ihdu4PsE0ZoYrCEz6FThka4mY/SZnbYXY8tXUlqOONVYIc4qf/Pw0PRqitIIwHeYwKyXHlYCWc
06gh/Q/S9uqmiOIjliyxtgRYEHoi2rJUhpN4ZWdcvi4BWI4VaLQM8FGe6u0nXg9l4LMpnM1x1lyU
6St4dJcHZpP2tSrWGY2mvLseehEixh27pHfCAW1OChJuJGm8lzCrqLRl/7ovl+w7O/DuiEwIt7lI
YAxtOpaaD+A+1uLFwLKwhE2iSUan3llK06NqN4bZHxPY9PzbaEu3mNdBS77CvqE1qydVYX5ttsZe
y8M4qBAeHExp/KOxOAC65ukrfppu6nEBKu/WEThj6FIj9yx6Z0Lo3O6i+/TBGoaRK5DSCbH9VQcM
2hkL1XUoetEi5WH7Pm44fjZH1CDdr90qpc3DEY8+4C1l/PjOBKJNmKWdIGWopezzWYm6DcCYJwFA
+KvwBipRqn/Bvp3oVXYnkRMM0j34wXV8MHDWpM5tSJKSnBoCbdJK56bwPUWhYP/0N9rH4JT5nq4V
8O/vwRTNR0cFVFc0eS0YhyBhG2/77L4R4wI13kekc4+T4+3vInknODljZe9rzXn+bkr348v3onYO
w/6k7DXl9tpZx2tpEeJAl5v34BJSmHAx09hxDxsK0996lWGetTL68h+dl/nSCAeSOXq2rsS5pl2C
eyU/ZWUV2hPr2Mc7gpKwA7QyYq9Yhk6WYHLELWpMxmDtJPBHThbNCy3oS8QuPJ/SO1EORYsoN7oq
dLjYRnKTF4ecOtHfKGDVc6buyDngj4GJ/OtWeiSwzW1eFSwlNjKF/6TCgHVr28TmWTLiKhv2pRr6
n8HnRRxngpq/6uKyOiSS6fDAluzaAwSR8C9+2B37y0gYpJYi9i1YN2peIMNA6WpIPiGwYDtUvzVb
0BbUn5rSonNMupuGNR2wtG+swQ4fJnOTkukCNrbtg0R9ShBC0nyIHwaC1wB7LLJgYpT2GippTU0g
UqIcHALI+hCJJTxMTutqBDzSmdpRrfW60QcQk/hk5lLkeYM0KVSobLmN9zU4N+W/eUdawY3nhDSQ
SGCQViaOI8LNqS2I+aTVqp71adBJWW1HtUJsMYUFh7vamggxWW3w4TKULcGWVGAgU9h9p4da7tQa
Ermrlhq0OsjfqcqH40IR8Sk0BL3dnz9om8DxtkN51z/DQA/pTk5lA77AJmg5TgtANkv1B80WS0Hv
rfhHg2cEXdcstMtlRqPXpg4L4klqoltijgibE08EAXiZS5gvdiUrD0paibAtBxMcbUfkSYzAH+X7
FAcCa6tAWP173sPaEerSCVmzwQ1w8OsdJeuWZG2s7V1m/RtpC1AQZmr/mcu+e2YVOJ5LZf2ZcvKp
GMWsYHt1AGInif8v/QdwQnr2kkUfmONlCk9xLh7PG9xbpPvW6GOeNz7HZZuK/f6QKxm3yNI/83eo
lzMbDTSdNgUabTBBPlvtmKAStGy0xjg2UFd4g20/EasoZKOJ9MQ/C06Ms3Df46Y9l6yylCFm0YG3
+aIhpGKtnv9xYnhhppSllAgRv9GHNKjFCcFVixyrZlHfV2xU8YHzsVgm/HIfaoi6c0+uMZLolUtE
F8qUsRwxmwdkpr9zCnDuM37f543JtlyZ/r3xZE3zBs95YzLjeGWYiouhhcOb3fOV6n6jqOFJAAlJ
yRXQ+afcGtKCcXB1FrWTsTFicwnif7SuYTrgBPG3TS6rcPzorHHE06059TFezhW+/8KIuSRwXgfh
26CvEHMO9AZlpZkcETssnaiCmk38y3P5iCo3OZp7fadQNcZ20VyK1zoYfTuClKS7NKKYT4VXPYOU
kK3xj649C2bV1JR73MPyB0Ov/bC94JVhF/E5c42iYJ2z66SW7ltS+jOIGlqrXNhQ9DJeN2Bcjkjl
SgikS63+5Nlo7+ONwMY/Vhwl3V9iCgk0NfhT7JwGjyRUpJKZy8BdnN3hvM8nEA/gWTECEgdHAZan
rL68Sfq8+kDPBCZHyWIjotegQqwNIWpuBprGMfSbSm335Ac997sKx9dBQ37DafhlWH3PZQuvT6wt
EIJ4/m6h83S7q0fAUvf5zAF/bMqeg3yjvmTRBXl7iwJLs9oPeyvnuwqcvEmf5RPObLEVGMV75W8W
dCBXm2Gtayt2x4ruvJ7sHhBRESexxiKdGz6rT8v+J4V5s2mnMFVcAz4yKmcBE0FlwSZmIfwTpAQ9
lr/u/iUpQGWrX5fyGmnEa/BalUjsemmwfu3sCvf56ONIocGX7NVk6tfNJNVM+8UNY3DhLPa9jbmv
VYHXxEJCdvQWLeJLeX0u1FLJaYj8ocG+hBavDlu+EdvGhhHX1pLSbw6gwxbwWAeXWVgFPXHTVPag
yagkt9hY2No4pXC7nB3yKezAUIUR3WLwSVHCalqkdJ2myJ6tzW4eng9kadXlcWjzdwuT8eNSV+L8
d6elGpDIETEPjNXoSaV4MSsEjl0o3gc/BQUkclef2lxRHkTPnkbbFD7NBc8Enn4GYjAS6a7HY5tt
cZH55zCLX7cyG0+8b+aLn/gOboLC49GpNkpk2wLa5BsMR2quxkIYqZD98MYoKh6Y+pDs71ZpY7eB
ZIM/r2xoI6aY5s4rwuKqJbAtOpzft4pOvCCoOOhccPtVZ9iK2N+ip7WcHcVt8YndEwAq/RbcEpfv
QA3vNFvMG7fcBrDU9tjULxxxU4NWpsWnyJ7Kz+b+Quv4pvh/7rqTrQrsHWvC0w0xB4k519A6c1F2
GC9IR4w7jAJuu6wv7sbzdvfuRtsHsGFXhznuaDK4IuFzxoxN7chYfQf2+JdZCLig51OTduzCs01L
vv5XSo4RE/qbxWvYTcRf8420oyIuGsCp9s1mn7enD8bWSACwRFj5/vMLQYfGIG5PjdxFfzjSSv7x
m77uV961BAxNUyk4zZJ+mpmbJyag4UiL0EDc1fXb8Pg/M3I0vQ3rASdvqkR7tG+oZgj5nHMSg79z
j6xTWW9yvoR4AZiw1/gog2Xsxj2FeIZ9utsAYeCSNB8teJA/4ksKC+QA8kIAOYUYXRN30ap8HWAf
2FiAbzH6Bi991IJef29y9v/yU1pwbpkrVwI8eGvs/apT90UbrG+QD5DIKUPgdIoi3nI0W901k4oE
F1Y5x/uDmUwuCZZ971rSBhs5vxfYBRjHStxqa2yDmDFumCbsFrkdxkGGFWUp9Q1HmSldj5OVsKMl
DdS+z4W2wvFb8jLMR+KWh2+yDEtSBI2P/Zo8VygWwtkwxdnZ3n/hA1KyIWljiX0YoKkDOUUv1RtE
mpczgcwHtMucY+IQkRw3fsr5Gn9gObwErSi9XUWm0Fx5kT9WrOjCk3x1u+GWoJEcvIdpEagYFLj0
oYqHOAqv6nqPDnPzVgv2EAzb3zDvFQ2qMb8w5RjuxuXVJNEMCSLZseotD6hDShdCX0Oqb2i5C9oq
sHy/RU0pnL+ofPiYUTMxU1GCr4qO3aWaJz6OK1oOQ29/FD9ws0vVuat+Bl9HBY+jf+imQU1VVWc+
1u88nY0Mg0U2fAY9TmhCMFjztv6Cc5gwtqoXR26Yt17vK5pNMfaDZSb1QpGggU29aBP2VFqjwnHA
j06noo+wltvuQ7mgJ19cKuDCddpN9mJTOX3KQ/R381NJvID6TNzLkyP7Xbb9OUjG6v1MaBcnbFdl
zo+Nu48Xom5n7lG9hyH5KEi2e2wV3B9bHdHxDeoalqrmVIrwFjeQfuVKDJzIX77lT7js3D2jVERh
1zXj32pVTjGdb58dz6I4a/Dl3XfSZRTQJ+sHiCSXJTI/uNtQMbZzB4pm1iFiXTXATEmi6mFoBoLz
QR6xYTry/fbNepWEdyFgVta8Cyogp+QEYb8N8uSBfRh8XHir4Zw0FYIgzwVDB4vJn81HrVkklfac
FuQAtD/rImMGTs4yRjKISz/7mbSk+Re5DlUV4/hpTdlBIarKoPDctvrTVmw9AZ9jA5bLEjEHUOR6
tXbeu9juEvBwAAk0vS7aknw034pslBUksp1GIMgI93zWS+XiYoRsqLo/TVviFSRN5aRicOqFds58
lqkhmMwikY/2aC1icTyIUvz5vB2PJQ0DDSskYqeAYx0mcFyWtP234b/B7Qdr7tIXAdpKqN5zZlgi
SMwIffjz9j9Rq7ZTZWX2xnKI+3p3cSmkOqM80ACqRFF1W2mOFnCC0vp1zL1NgSvzACD6owfjB/eu
8LuqysKrccVToO3DWPX2YtC0St7Yhpf/3BiwfhmvrKRByyO+iSZlbRSNGRg0O+TC6kMvrN2R12w/
c+bRMElFzBfXZo81X+1zZGzqBZMrHsHS86+CxbpXTXGgP1blaRm8lcpPiDIkYsA7s6VunyAuQGOe
6/g3KTnGaV8HHWe5JnfYDa+WLMmKI19wJzMqaB3o2lkOSwZMujR5LwjLRGhwyYOwKdEdIEht+7ZG
KoSpMcGaAq2hUbWnQ9eq8rdIO/jZUMfwWYtYq9sHKjteGjFPeG7I1TCy/vKAArlSaf2je2G09PAC
tfu0z1pNsqc7kdoTMs18Jn7on9iIjc/U/MELYJ3X14CpQDXPUpnmHOMcRl7KRQDTf4oYzGqENUbG
DDCDT1bjOMYTmZVS9MisPzp8pJdqDlBKAgMMC9vAUqR8FsUF5U5vKDyf169hjbDgN7cqAQW20YSJ
KF+Ob3ROiparMUap4IW4/9/1WtbMCJ9tNmUNWqI9bxnrXmYEndxK7f1ALYGDb0i0oEpWmktGyK9k
dEA4bVcOV5+oS5ZCtYaz+AlviwjjTtfjidyLYSHrX7IWQs7TfEmhNgCSr6PCnnC2nBu6esFl6w1h
9Djsf7Tti2Ejr8nAla0dLfZBy2rT2yjfkjAat7CJITUFavXcDCorQZVIDsQYupj0zp8Oo0BKBsO3
YgMVjmc+MjAlnffY/0rqPnJQlDeUbRQADfIQYFRs98QRqmJHbwmUssUE6J5kySnan800+jC23gcj
f6DFxgW4+U99AoxBfxHQfv9v1qmTWPiQ0neXCSFyV1jGN/litteA2y0XbfRAk8O4tHf+AasAsOhC
UkPCHCeCzy7DPDtl4cnQldS6PIVadiLSnEGq30nxGCY7ve370pxFl02gck3kZrnEdzmRY+4PmINN
o/qT5c3nroAJWZI1rKyjsxnGXHHuLfCtz3hThMZyJV9wjEc266zqEBnZXVd7tkg82WwByo9OnvAz
iHzwKYOJkuLOE10XoVFxI6MdjA06cAhCt2QrdR/llcmG7aYy0EEQA92xNDiMc6nwg0HETdwmxLXo
1ZvP66P2rginJ5CQrpgZv6ZNjTYUvpCLRbnSoUkykdW8ZCt7JH+TA+XQdLNUSnA24c1cejvqLLCv
4XpKQv6/APMEpXOYtBgcZpIZgH7i7Iqyfhwn6OmX5q7z54UU9PFEAoCZMQhpB2WYhrsVOnDRdKIq
pcmybistLFHSX53tLYUVqJMEvoEMwQIp6sMVpL7QlUh/5teqYZNMWbly21+c11XngCLXc90tiAYk
Lv+mmSA3BXjcmUlkKnHOZjIL7FIpZuUiIwcCfWKulpTFH4qF9LHpAVA2aCv/LFT5N5G9M6xO77On
unVPbWNNNzEZ0AWN1jdtkkq1787eUG+crNYQABo2k3+irwvSIOdOcy6wXXdV+Gb0epnTI9nwXkBV
0ym5d8/HQIOp2otsAvpdKp1lql8/VnpcUvLWfAUSDsEOg29ENefiqYHHSgCHDquNhjO1WYwQvg7v
VIyfuDspLRY/oKKIT0b49gfp2Mcvd0Uqs5vI/N1GrmO9wqCwI2jV43rTlgop8ESCz12i4ktKCd/d
0oXhghh+DLN+Jsj1hD9QBH45kcecof1/bTb4sgq82Hd9bl5wE8yxdGgXf+BOkncMXptfogLCjAIp
n65iU4LhCQFD0FzzKlm87dL94a6+h2z409itBJa1rGCLv/NS/DAHuSUQfhBT4p4bq5ftNEH+ev72
nO3Hd1nakVAuv+Let26cLAyPovhLni/q+xg+yR+bxxV6ekhwr/vrFMadJGrcj9yNQMQhwGxsU+KI
QKTs9rX+H0MgL4X6mZXU/xNLlhUoIC8RivvH/yncVtS0yaIbClJ8YbnG5AtxWcRr9BvcGxaabKyI
59zI+TdMAzmuFm0A7sIcfvhPTOLULAwe9EcPLbj7Xwb/x5Sko3bt/DFdga0KP7ElhuIkP3uXC9+b
yU3DkCipBA+nC8dNW1PGSDaCCS2MZ05R9ic8QtfP9PPjtQT4P1NxBFL2w+lRO5S1/UfGdqJz2Swl
ld88MQjEtvpDmFlxxCGOk20B+DkxSFrqzdT1bzRgV1MmlmC43saGqy0JFQW3A7w+XzjLdI2H7VPm
1VgFyzMevD4hblBJaDYdcuetL583fQsyFEu0hOE5gKnVhX5oSNzBZiVsh+cZ5W9GP0Zv3rJKeUA3
k7YhAsmeqziNoTEfpyeTywrOQoYxtK1r3cgXW2Hj4ad6TU1K46FsVaLWkP18ZsN8PMlE+6q2UFrJ
orW7U0Ba+33ZqFNozmWqmzAd9c1V+U77UtIHthjQnWGvCc+08RxjyJJsydJWuBFzjxZ3AS8KtfC2
QEN7xyZBLGH1vrtywYJFVq9Jt2T8r0/eMS2m/rEFEvic7ST8lg1pUnVGFBwsNuXuPWQPwY9kU6G/
Ao+TrWJkE2oetelrXPVi7+f4kA5lHMa2V6W45qauroslDu80b7wxwzZxZWwUkR8fmZ98AsFwO2gb
VsIeB/9oTbBdpleTreSFEJ7VwnizuAiYwwb7Kh3rlfLBjNPOomdYEBGF2dY2vHREFA0eeCHVAEDh
aowV5Js2q1MkELicS0M6/4G4XjHFz+kXaGdtv5Lj3s7bGHnCjeVyju2MmEeZj7KwZjlU2vcv0NVS
sgV1VpF9YV0ilF4CznJN+wBGpjpO3z155wRDSTFLyOReAYDxZK6m5wYG2kHDDSf0PPR82ME69gIN
AfXdV8lMh/jOEVfOn0yDXYhEKe85XnoNnsw5d8sF2xJKNnia9IbsL+NcP+LbdEGAkZEVPMf11d8R
5XA2Hv5iaflqinD1yL3aEKFlftZaL4Ph/ECQNUK2bhRdH187uFUSYmwyu7fKixXi3Nk5FkCULpsw
r0raXhwiEjjCNWrU0ETL9CxoUAd/k8FjZ+4JaKJHGu4L8wHy17lVcK1ob+JfsWHPM9NZphJrbofg
e3pF110X280y5u+CxJAa7o0VovnCd6ijLynlf7q2a9anGVMwMkmFSLhPkSnIDOiDtubmw9QEKeEG
xK0V4ZEQiLhJcItVvsjBWLQLt/FCGt+gV9Zawf2KGmsktzdTa2DmpqOFtTmNA0rrK7oFnID51udl
wcwStY5DF/pwXrS3Sswts4gwrQINOUX98totvWCZflJQ3XbQh47P8zPZDryAZvQCecSIwD9gERvh
ChxdKHZwSBApGnKMvL4rHHbGkADGyy5iQyVrUoF5xGDeTdKkDIXKQhT2LZ0ZPuZ85DhgETr+A57i
1fWydNjs8yQuxrIp34CAB2Q4clOpD3TVoNBTNHc9bk7uo/HFmiJEW2jY123GzoE24T1PgNCkPARn
dPuoWUy/V9Lsmp5/VAuL5+4r8gWoINI70/+dXSU0k3yy6oCxy9HX9DFOuWjKYB75+0U6hRNWZZ/v
mbsdoLqluTAsS8byBdltjIcKeRX9mDd7UwPd/urDcXqW3guvSRP6QvY2YlodgtZzy6B38LqsTQO+
O9d49nQmJ5kKBQsbcq9qijto2kk7Mf/W+1k+zhncKpiIX6PeihlwBDpetbu9v7dHST5JwcEhHNqE
U1V4CZiUqF2mW38PbvzB4bd+c5BDxAF9uwNPTsmJf1aPlci8L5a+7C2lEPADdSs+OANqyCqurWke
YziddtQVz5S7PB6dEawW019TSbQrgbPDGW+foyrbzGwKObqInFXuzdua6Ja+N+qGSFS7TJ6XzznQ
TsgR1LLPsWnlst5h0CEsA2oOSyRwGbq3hu+dEOBZcL8wiVSCNWnsHjf2RqU20k56JQ0jwP4aK9/F
EIGQj+c9WLVvfh6PATzi9GmHqkCdZyzb8gby6GKEsTFSWtBPXpChAUEf3JriG/sdkh8fG7BCT+KH
Eo984y6tv9eSUEpI5SytsXZjlXS5TGb+oQRWDT5EM07cgG779C9kGpf2wO8z0PnyJvorKpnuEbqp
g9HlJS7rN/xR+rmWurrEWwud1yb189R6BHoEAu2TKkGtmoYZI4pClSnHfzmSr2gUXMM5AYFlT1vv
kLDCABD6IrMUOrGbx70yYP8s4gbUGGtNIZkQPuad6mZ3mtIRuz4KYUwszsxlFYIJUzWonrtHHbVW
3GBsuyVERna40edOhEuxZfn54NKCfg9KdJ9RFp9dnIVZ06zCymzPWalKhCt6abvQ08S8DcTl5pFt
T826W85p1B3Nj9bIvOZWFpaYcX4qGlqSJpquoywjXjs38HgEnm19EnlNWIS9IPv/Gcr3Mfz7A2Vl
iFVRg083+ik/kJ+kuYWwT7ml8KnRCmIZ+WSUwJ2ncYurUXHCxK0TmYg8Zp/58I67i3S1rNXB989K
UifFjsvWYktb4M5SWZdaSb4bq17hZ1LLMaH/In/S17Z7hcGx2ZeFaksGUBngV2OiWg3IzewEjyBh
7TNSWkfszdEabqi2JtbcHLupQLXZ5yZdPPioAMZIOHb8WUFpjjY9usotqDleXggCajNxt+2e/xZJ
1LQorthg8lsZ7Lv9OBICQtP3qDg6+umOqHT1vk77ZAocE341wFKgkkbxhks/aRlmoRGNwb2vkI1l
Ws8vi3mEEINS51AbfdEecj/zNyjL201faCM1OV7cbKnfPQbKYkrRj5HsWZtMRZWrW91XZ2FXig5K
JgzLHhU9atPuTnQ/nofS9WTxb/x0+2/QnBE9m1WYZOKSjOFqF590+qXNkxIU5aSRkZofs1M6IrWw
EamRr6mfo5aSelE/cKTe7cUaBAQW1flMPgtCS3KjhTyArxTyAnr2aExNWoBkVHY0LxDnVhFNjMf2
dwo57afhz9mc7TVn9p+a0M/mRqy/uT/55Zyq7N7wu5QivBN/J6e/fcLcXWaJUf0QBU219R3OXnA+
vb+yAZLycXM4Sb7n7C05FM51z3S7P4mtV2PQGqUojp3ahCzeX9MnaamOYeNNjfsLZymUKXc+nJxo
2pjVfMIBJsYW5vR5KU+Rs93fGViTPpcZ13bEkPPpORnvaOhEjWHaNGHTzqpQva4gSYuyhxTFzOWG
gZ0VUFkhDhuRuw85U2ikW3X/vvZ4Bxef+0w25jVq5daTznPKGhrP5FNtVVl+I7gqbuA7L9p9+M7k
dySNDm0nhG9UBBu7g4AvOVNr8u5Uj/WZvKProONSNRbk03iNezTBjtZME6W1T5nwjJTyWai7HWK1
RwTeROhVgm2BgI2Re6NqQIBXCbwnaYdFqjdRybKuO/Jd9jiqInXP4EWZfNGCLvVtTBDO9WR2glda
awh9hsftzU3eshXfnMdffJxEJ/xGmSpgSgJ55gNJvgoL8gWdSb1pLEFnBWuCcXwEEoa6JBo1a2+t
u0xKFylNMRuhhAfka2J+ltOhOmZ7pzBDavUg/Ae6R/taIUARKiwJ939J9hzsykN8weXmz8RMzhzv
tKARft8rzXwGqyXjg7sZXhvZMN0Obohilba8582/T2BE0D83Zg+M6YI6BlzUuKLr/Bx55LGocCKQ
M41XvaKqP2S2l9nfoxggladHh3uGS8EfmlODONxEkYDa4NdnIXnV+Ic49QfRNN/096d0kdC1dSh6
OyVPggjyumPNwsV8k1p8qhbFf1xyw1y2EdZ/juvvOhQgx7UA8lD3YG4JPbZEFrTeE2t794nOftfI
x5Y7n09rjpEHzwUTniY+NQGSEIqjhKGvWNYuABcCNa/Z6+uAw4LDXtcoYarfgYv6CmfWuMRWDchq
9qigohZ+NrnHwTuJXNHez/LmlNDKWabkT1OPo1NGNeHGnqulxuatKTPF2HcOb2aE3wIsMY3AFaJw
eDSnEj6SbfMVLzaxMmSkSk8rNzBQJ7CcRoWAOicc7Q6h8FwDlV0rRzRzVpOIFCX3Iax2WQit6fhe
ivVxV1K63r9XYCJleoeFQ+bgqfY19oXFWi9eYWdlZm4J30p6fVNN5VuQUTuuHhAaG/ha1uKiFQt0
0o8FpxSgB8zfdJfWuplN5dnf8ICSYPDXrtqHtFffkXqfg3TGBIbIYKNbYOssZEP9mHegbylPJ3ZO
S3ja4MoklAHZ5VCagt7tbIXxvxDrtSljxVqd/887g1vJJ1AQ2uDwyKYqMywOOYuYW73C54DobYQk
Vs7EWO/tZ4/CaFSnvRYQQYvWLaYAMOelALvh5pd58957CUPRJ/xYtVz3e+UwAgkMbfRDFn4MQ2vs
iYkgFD5hExUziPhMRXSURA36KRBX9izHzbQkyvEYplGatpxdpZT9rUtUOZOZee/qEGEkGb3zSzUn
V/TZ7oXavNKWVc/49eoSTZm5tAKhenI5gmEAUsWVPvDyGETEy0XuAUJKYTyL1E7CWWcn7Yxa94Wh
BzRB66gLkzGIHKXDy3fFppSLJLpnoG+mkKdFvpMytl/T40GQtrUj5XxjZ45HmFxipGnebiorSprx
N4m6TnkJqAm832BeNC0t71lH3ibtBgTek5D1gxWojpNsNpcmCAjfLuQv/XKeHE2kfJ/EiN+uLrQG
Xx0ClCVee3jdvW+4iiyRLKt3KJkUZ/uD+kZ6uIMBTmSTAMCxk2hQ3zjZ+0CVrr46sLTjxvZb5xB7
P2L88eCzWV87bG3eWnL+09O5IXK7Fhzjk1ZMKp9alHT7qpM4spIUdXIvFEhppEjW4Jm8fG23461N
2ZDCMh6CCh02Asf1w8CaKBnreqiZ9Mt7p9JYqQLtEs5Gb5qN5Usa8PmPZ3pFsjjPw+mY1qy6kl6y
BpIYd5ymPxsYJt+kx+eL3qE43M4QPCWJ+IzhJ5L4obH4o5D+3Gjl32Zjp4wfsDZ3z+tJyzZijHdO
BGSaISk0DUM9TxKtWNo7FJ/FnNOh9HmbZaQ0b70fMr7MORO4of46MZQ2TJIXNpqe5hFzJ7E4d6+X
9s1CT1eUb6jPFiJumRFECnXTyvG5kDWuCi/+c+t2cpM0nA3kHubv9FiYmbGxMPXZ1aPQMuetxkpI
YLDQoavgdth9k5y2RRevEQnbi1JiRN127x43y4qhGKerEqS3Kt8E3Navul0wv6BMcDugn4x9pSzm
EUufUrfAJcH/lzxupmbU5KMS1UNvG/aNPL/yB26S0ZU02tSpjoDFFBZbq7UbIGBoCE2iBJ5iwogb
5aVa7QLxqAhPqhKB29yzisavsqp28J2oWrFNzbGEG7JvluYzSdMQ2G3LlDGvHhtiSrJ8QbzRsp4Q
boysZkFOH7VztKs22oaN0E3oaV7JgqKOn29R/33dFRNvDVprGkd5kih6W7uqgIYkq5JwNWh7hbpW
9LGunisqiSPXF8lAjNrScD8vJrUc09kToLsSCC9mFiefuhTLrhX1SiWBhpW9kEDq/AfMHFiVZ4o+
3svCsvfMDYeuZkH7zr3hYapsEuf3Pf22yWldTfLpnXLOon0deTZe4azF9s1Dmqcw8mCXZX9JHYyl
40fWegOC0Y08GTCRmSFDHicDHf/HkGOR+p/DIMwp91JFeE+y/RJfw9UezFuTFDxk3azAfHPkoB1A
IyD4fUtMAJByfpJJayL6NANs9G37n/4foty22Se6LIXSGERy1/RrCiTiHKlBqjGXpz2fSlde8XR0
WLfUtp7mevNak6wnjucwzlfckizlqAJLM/bOryCI10aLoniRv8oZIAXOKf1uVG0K7CuP9ltoNxpZ
uMK96+fXdKnlQa9nOX8XAFVFYoruH9Xpqx01Gs/X9rAx9XiWomBRIfuUpjiAZV2ZkGCTUDMAw4F2
Iv5LDZdoPHA4/Dj33SuB282aQ6wuWzgiHspxMw1H0RtqAV0lI7H8S6fPeWqZixrS8luW2SeNlmJW
FKSMGuicnBavbfElnvhy0x2Q5fj3Kf1DJHpZY1txmZZBEbqOEwV8P1+rADqM3EgWsSKjfoR20e51
vw8ZTolYhm4VmZTrF4X0jBi3dGdgKkwZySYodJ2dxsLlu2qmAXjbjaUOgzjmPS+ZLg6X87MpQHhW
dwYo22147aBijGj7OqK/is9buGP7wjLNQr+mKnAU/SF5qj9fNjkAyP8RuEEEjgxtQlfeUDejZzz0
Zts5LFAICehdZEIteKfjJXyY12qPOEWz4KlPhvwyprp1rF4RjTYFl2bkCQMLNt8EXqn+Gf8BOx/4
qDxcASjugJO4AtlgKsyk4WyoiE00E88vZVLPg2IBYqSfECFJx0wWR7hdCMFfqZrI3WuTtl2wAYZJ
gwoBblpS+S8UrdCv1JWETJ2KPyvS+uHSu1R55bsiAYoQokb83naFKA+j2cXm95W7A9FuLCdFScLi
4EwHUYDdjlqIKWjFX17qUL7KWtxkKZKZEW9kM13tGqgDexm1uOPghuGfnNcUsHfeDfShvI/L4TZf
YvPATvYxEzhNWvSqx2kcZhOAgoJ05z4mg9sJm2H8e3ys59lWqT1LVe0yLqNZAdPyjEWsMZq4BkAv
RRbAG9WLmZDwhcu81/GMNF0Wrhq/HjimRDYgl2EzbGfzZmN7cSXePdqA6wd9kYz2lZyeGOCsACKN
CDj3as9STG6cKfszTR95wGrHkTE1UNIcDWOVtIXqtjRfqF71dxx0SVR0imzdG10e03+DfY6zZwhk
+bCu/LV5RdSskShoTwAdKmfcX36jVYTmMPevJeQP1zSzkdPghOMGn6nqxIdsvKS3oZj8Qi7nXiOS
RGU2Ik6ubb1LALxhdfVny9Zo6R/SBCoIlFuWXp2IHB7vxXOqzlb33x0D3odsjyp08pDpDkM0s1cc
jYywrIXcRBWq8otewW+jPGufAxBYLK3sHt+GJZ6DEnHnbWIMB23EiiLgVp7rgHZN06Mx/2f25Acd
KUiRuFZ62mhvi24w5cYlReD4q++5zNBYlvLijnU3VDH9TzApTfqoBH4fpkyJ0okKs0J+sY76wi9S
i5YC+yJ9+mIKrC9dyKZR4C5a8hxRnzwfCnwvsv+2bSAI80YV4iKJhCkwLBd4W8rFgjd+l72Mx4OE
yQi1BXVCN8+wgFIB1JuYQZA++smJbySxHabVAPBPn5/iCzuLROklCYyx45VUhqzcDzGPUTeyLKuZ
M88xY1xcclVeGnxvdxknQJ/QaP/95flsKke12rcpKFWt6th4Zy8IfrTufcjE0nHIBIjZ0wJsJ4Ho
I5RVKr3P1lZuaLTR5Eqhr/Fwpw9odDyeiaFePc7rkbCraQ6es0ewCt05GMbi/6/x4o/GVGm/FNk5
QO6EI2X6d7lZdM9L4mit9a3jUvVSPDtY1JKIcKPMsizbyZlz3amt8mDWDK4/K4Lnm3YnlPGHJT7r
FHra74l9SexWvSKci/nM5o5Gk30Tk7IqQFeYZO1sTN8iHMCQfHOPGWETtYpMrGsl+BTsI8c5Hf/A
DsrJ04X6eeWm/I4oi9pms/sIPXVTqrlJFE6gjxu5xgth3AtzD/3HZLiBOlTFORDw2v1fh1cimMwP
XW+qi1f+1zpK262EJdIl9knvmu8YPjC4EEiEW4/kEUtZyCMCGT/C4Tzn2K99AWKajN4hPoEdC7sH
MD8n7/PucdS2WRbMQRBNA1Ap59cjnqHU3W2M9IU4AVO/sPtycIjs/LzbKaMdx2iGZeKe088srf3C
l9w5bbQ4va+tBslgfFf1UMUExfZDNN0Aij7GeglP5QNVCMAx6e/cw0uSwg5tjQ4z6oTEnk1hZkYw
IfdNwBg9rIbU2dGivANE9CaKJ2iAg0qrvY+bD7m0SZWrL2nwJB0ExyQh2BwhkQdMa9Lwc8nRDgvu
SqwO8NRQa1G/SkBvCaiQD0AJn1MOZN1TXpNbjpyY24V2eE5a8RAaWG3cdPPFyGZddH2UVXYc6tQI
7VhN6FctQGO71n0Ug8E3MHsfugCfE5eIAvDwpfNBlxGqOceIoAk2lQd4tNa9BrerhiIoEnCGB/nT
n+POSEQsKEH/5dcKvH5oWUdBKZpAcVoleFatItOKr0ExLK3bP5USCzy/AWuNA4vn/B66ALP0Pt78
hYYsNZBwYTGhHQX2S2Pd1zxE5hfXHHsrnrTLUvA4VNCkWXj0Ten1Z/Z3UtN5m0arDCcaAl+EeKNZ
k+MhHtZOr5b8enq4TA3RjrIhF8oQOd9PFdDUK7usNXxPqIKzTjGOFdzo1Ccg/s7lbg6SfBpCnKyO
/frS+acRs/9ELrFZJZghuanO8/8vKGx9SrKmPnBWmrvv9AorLhDBYCbP7c8YApWYWxfyGsygZ3mw
k0C+MkfGYgdR9j0UVv/yH45rpvwVmoarB6FiGKXNx37Boe8yeNBhOlJUE86gq/z1yb6tbNSfiZor
PPeka5wMKJau+3AMQ0CgrskWZrJ4G8Wod+woXVfQCYT0BVpU/CEKI94JugqHlFfRBiob8YTe/e0F
fLuX3Ug1qd26zqimfN8zquZ6rKQw7/wmF0HrOEEJC37YRYtsh8BZO25ZsaRpCqKbhD22nq8b3GJC
Ehh/ikh4DDXNehzzleFewVqLNf+RVYntRw3a018jJriFaBQQU2LCkCUaw6R0zAwCTnvgXJnEOvxT
rW9uQil9poNWIdK+Z8wP92ZljO/c/dFA3q9TbBvdqieMdtgggzSS8KMGyjoIVFOYCeo2aUbNlhm7
XI4OdZM8P2ORYE6UuNfqI754fNtZq9WZe5avs/vBfIzdJcefH0RKhlp3gCu5Iloo1SReH52wmEPS
ZZum6buHt9lkaYr5/ZV0EkxNfT5R1h+q1WeIOMAMlCyRrKHgF1CNILTf4shX8FagLgE03AVvD59C
DgHiR8FWWEQNW7wEXxZ89fXWGWZEWLwrmptT+2zG4mQ5DfCgdbY+//1DGCjoWnedKmdXWaW7ooxn
OZt0s9Na7Mcfwj/491XVIgyGz4WzG63dZum1DgWNNv61aB38Hd7z40Rp3RxvfkLuO2QxLatktcQR
pNl5Gs9HtC/DHPSnkAm0SXl7Ld28aP41srnXAOCG8cusRwX47jYHMtIbAnZcWTVSTrTtttmy520L
KBaFk/DbCKGrWxDY2u/8HpnWxt9BzxE9aRQ22DTCSTRmuxhQfVMWBCiiFYRZESK+0tscW9LWdVWI
9ZcJ2UH2F8bPMH1b5JTjC0bhazANx+liRZdCsOUgXrpcMT1jhPA8OznnqKFMvdsZorJCknXKSIO/
nqI6APU4SLhSvN+HPIOy7haaXzoccDujnHbykDdqE5gJoZo5P4ZW7raeoy2k66BY1XVvRrSqGGIY
P1mcVvckOUxp9NZF7b4UvynuOu4BQ9K8ytW2iBSXItjgpzsAYkTmAmOinIdIXkzI8E7XhRPfPp9G
D/mOoQ8Sorgw7WGu4F+ik0w8OJ+ZF4Rf56hjGXo/mu/AvRN84ueBLdRiCzFR3GeOOl33IBdFJ68P
iFCKzy1MIsNMRizwYCP6NlBj/ybfiYPdMsHTYc7x6rptidQNxjkCjshRe6eBR8MPzxnDTS2wz7IF
njXbWK39aKt3soCCXYqFSUyyQkOZQkJFXmdqjiz5MKR3lYCXpZ89/fy0i1lF0EnMogJRCG8adW5D
Gu/TZbq1m0G1WE60bEFgh8nhLuKcBXeIXsxyJJa0pXy543bqkMVd0YDZjrfwsOeqst9XPefJdh3n
L2+oz44exUunrJpJSaPvs6xQ5cdbifQBxkIw9/iEW+t9RXOxa8qzSyY91pVFTWRiYtva1bKgkhhf
PAhtSKf5aMcxk6ZHAwvi4UPBRkktxygeo6/3QerLlmV5THpMHo3FWfu8sbf3liLLWbtW0CqGcHbz
ocvYH74z1GWSbHoBE63mcQDCpw8xB0dmVmZqVw53VmdwGkMn5e86Em5nVx9ZOve+jHzdQHIPUTbB
xCiSi34knZP7/p205qh62QHS1fu45NiGgqUH+9pitXU4WK+zeDBCWvFc5sm3tcBb/WJFyxH0XKl9
JWRok8uMeUTeh2H1eWUo9FI1kfT0v/VWgE9xCcEJfXtkUfJUEDqjOc3/9s9IirDY8Fu2fnMFRJcV
Oan8zrjFvsKZxxF+lPtlrWbB5/z9P5Hgu47I5BNURHbDNuanK48gag76uXojMHTGIq2RpPY+O6pR
hSLCTxWGFDMnAg0YKW1Jv2omtuGN540Z3ptrAdb0wOF60/E4vK8ezgqoHunx3UpULeAFfdhNPVRW
KowWOtmmNhaZ/oC4eoggmCJsNBp8NAFkfO2Zc58DxL5lHbhli4V1SlkIUMDHdmRG8H0XlNOeXGwy
7mjV+hojILDK9fIX/pQa3duD8tx/9d7oa651gtj+UEoJ9HjWG9fJ9eJt54cdQOod9b/73GitlLAD
IlezhzBdzKgx08wh6nAAlmOfPScmsP1uvBm1MZ33ebv3dZ4UYnI4zHR/eEtBBpICshvyv5g/pPnY
cPClGOJ17ytdrEIrHS1X13BAWqiYmeKv8JJzLAn25eLHXI4lwHIe35pJoirLNKCupSfWvm5xisQa
eOY3e0p1snMCQwUIeND/czoIDTevWanvmh0+eFkWJOUGHtkSiOUM2MR4VWHRX9bJ93QEdCC4H6Fv
ManQnB5WXWcN2cyTaVSRb2GxSiwmbi4ik7KqtBkIf4+c25vugzks8YLoTxLYbL5SZO1ugKLYz3rj
EYb0f3/HsCJdMUb/onNokschaX8uDId1Sie5bQ10TfMygO2/o/mVvjc0LjgKRRA8vW2j2CKdbv6o
o9U6auOZYV3pqPxXrih+0IuMg8MT9IRmCP+i7GPCZF4i92GF/QVH1jcU2+eZWvi5pboCxOFz2EwY
b28Tg+fEzTTAmJRaNnxG6i95Svy9vzKzU5DGXX3zpHkfziaSr4hTY+RgJeCGjxwUlhlkoXFuqgW/
yuCbWXICOI0Tu79tHKTbHKbOIqNWtsVwN0XH/yJo/k6kXL1UsbnpTpe2N1I5MtFn9rvcMK+iFfB/
Nd0VR5/OpVlVZQwYpWdCKa4+xzYqQ7G8ukkD9UV3fZ5ZvlCaLROW7S5i0JUKjOSD9Wh2f/urX3KF
sdAYxCpKBhj/5vvEDh+kbi2ZH+TFjvSbaC9JubNxqc+e+hJkQgZ6CZNaL7o9E4/AE5kTRGEgQtIK
EChV772AS+j5dQKyK1jeeeN9zJDgFeVKNoScOjU9wLCbxR1R06lZEgsPa7NkSPeLt9gUUQXKB91e
fc1bWir8JgXTHe6BdYQ9a8nk+dzPVrlkH7WAIMTXzeNTAZ36SCNPN0cMa8q2l6VBEWV4vguw1QDL
yGjw98N2wR4773i7BuUo76NC5e9AenfHX9bzxu6rkr+7nYcsazbgRAt5hSZ9QncwFC6f71vvXuda
xH+odCARatv0S64/BARnHmyn5LV49qrQoThTtWahIzGdhmNYF20Exav0pO0xqbM1b6bjBDzpiLjY
RFHMrKSmOhoJxxm0T2BUq1F6KpPl0sWsN45rxDUIk3Mwc0wRd4i5wKfe2fV9TRJ0WnD47v294S8f
4HITFenVqncJOre/5WL7TvZXLawjHxTLBqxFIfAAg+oSb4J2xp8MISZ1Zc6fCUxVcghpjNWcQ1FQ
W4hBv3QmazDi7/2QvDefAJ7jjvOW/J02U03PcJfggWuu7p8fWuTqHjRvYf/L1J4zzEdYAxLGNM9Z
3qEBg7+uMOQZq/c1I4R8mlJyrgqsFByujWnLFddiQ6q4wxKYLtMBN/b/uyTDW6Y/CirwW+2uWNN6
ljqJzcyg5MHV419gyDxH1gR+84KizEgeGoZCYHd1QFGqa3gkThMvzjfwEBU0HOKTzhqOWuneuXIi
bBfFdakMKuQOaHyqTdyuS3C4YNBOCh+1MhEi2yxr81jt+QG6N3plPg3pI/ahXoG04PBUbsiMZOaY
goEtngshUAjQQEAOnlpKmhLfwZfO6Hp1YKtUiv1FEDdDlKk855lC115gYoktCeLtOYHmtk40K9uN
DimVjZ9dkFLJhqkBIVV3YRSINcNhGWL8UGEdc3EeX2ymkNihFiOLMpf+74RdTvb/H0REfp6stPjJ
1e+l+UiZtC0rZeSjdAGkBuMW4FhnBZQ3UMSGGxREASSEW4wX2yRLfZA4j9JmAQHUUT53ihL9YabA
maUNZIcEb94B7wmJsZFlRAyVnHsA5vy+hxgCmssLVVI+Fkyzk9W86gu814cTdkXxMEk6Ibajadwm
rb8u+OIqMP+65SWOLMqObV/jnDFiP5g5+oMEuSvXgeiJRugqiC1R3vG101SGhiqy+P+C+WG9uMt9
44dVRZOFOpbDmnt6nfpoLnckDebNet4waP2BNTZ/VSLs5Y7tJmeWwDqFLnPPtvMVwy7a8wd4q88c
DqX1OWxMwGCcqGnpAV9c2gvyfKnUhmMtVIOlmgF04jHA9l9Y1SH+gqHNEVKSLdGmNnU8w4+VJnHu
Mg+5AgwwWPcwYpAfQiAa8YBtG2V0JuS5iMb7zxXN65tFUhc4ro04LfXcsYDd6HX9u+FhCB10r49n
NRdBV/TMWq6wrXWYYYcei4FrcS8uJ76ZiG/nMdNpzLnVOntKvAdx5vVh7kvYax3MIJIsdDxFMcSX
WsJBJzHB6ByhWx2XP4aGUK/s3La4ANGUFguup0nTIkZfdmrcfhAicaJWb9VNmc6cBUAv02MhxK9d
CJYhjvoWMh9BX69ADUkLzOtIGiUoCvToBFw+z5rh7pq4QjXk9eYBTqMGdIpAVTJk+2tukGsGAra2
iO14zEUyReQsG+AV3HeG+Wfo757xvXMLvN3uoF3IQmo9RtpNbvdlsM7jQCCs2h+0+l2C1lON6u0e
TAlhNklv15n1xrdBhnXoQfdzdLJQel55k0vux/VOZOuBqHw2+eOOz9oM2l+xHW2egajJg2wqlnj2
uwKpvrA4sqQ6+lrq1KK84m76MRTn0auSCXJ3+Mt/UyrA5lV4Mw/PLBJ9OkvIAPMKtlvVY55OSb/O
ZFgD/ljsPQ1BPuT3vrHIoASOuf8SG9kcJJYdMAvL7IfWYmxDmBYlK8ZSXXHYOZ1y5zVtrzgVNxvw
LsegKhlJIT4kL7ipKlEvUwc6mnzxRUPj3hOFPPC984fskPPqG5YFlJKcemdzzF8/00+Ma7WWnjc7
NQ/FX4EUr0D8Gz1vHMIajcmMhPovsOiOTsj617+lpX/SVFjMqFFM/7QwPLlqNzywCTLQapWMekKh
giTjaYiSm1KxZHcxqE96/rIWnEkuby0KuG75rdfxQVyfvICifQyaQ23cg18gAr9S9AForzcSRbfR
gR1Nhnm2OR1ReuVBZRblufgGP9zokDpQxnsQHuPT/Tp5Cav23hvJnLxjG6Qfzju9DF8PjUbaDn+z
R1Cjhmu/CJG/eLelYYtxlyrxRjB8AjGq2nEAsbraOeOMmWzIJeV9Sjt7WgZWJ7z3jN3O+Q7UY3B8
vx1IUajxAFt5zBo9BbjntwaXOCeFeG/rwmgu/S0FKL8Qf4FkEd720mt3KQJJXM7+yl0kiW45qsVw
kN5JscdAtee+BcrZtYpWgaKcENRjVjiF5uPjr+zTHjC00JZoGeJ2jtPIWTWoLco3weg5gkEyUOw9
Jl5KmrNo1prA9WROiUK8jPD4BAEMqq4V+GRmOMc6XuXg77QEJL5TOoAVAWr2f0AktagyofZDZZiS
R+rEDs9aJhLY+Fmnj13jkcMrUJjKAfl0R+O48Jc6aFdYcTB6CEjKIqLgoER3VZYreDKrbbPKfn9Q
aRlE9olmR5fpQ4FViirnxt5m8tEObI5yflPA083oRodl1FX1TSnjLFxrdXFKUd7Oxtfdbq0iOMeq
kPSnfT+soag1UsV0L+zc+019x+xvwb+K+nGBOD5RyqyrMvS08P6+VWtq1rkz9as/WadNlFMG6u8+
Ud9U7eSO6m5bv0rTntILHfj33f0sl4F0rP2yx0kdbK6eDSOPhUozRjbM/As6H70f8AEcCbJRG324
SZ21fsQwnINl8wNQgkbCjY+Ghmi3OEccpE/WhRXQPmCDY/i+wwipm9Oc15LpRy9FkXSB2f9KMyMF
Gqt7jdBvi7KHWVrTTK79dXa5O3pjzN3E51xzFEW7Ge7HuUdxjK2hMg1oK8N0tieAwmBo6N9MxQDi
LnSG5JyA8yX3CwzafOKn04eQsoJ4uwMUNNfRlzvnz8nfGv/aKv6oBKhSItNITC0TKaOEKzvBlOxh
N/STMypurEzX2ZwufSlWFiBlAEZptMjUkUc8EfKtPNpVqigkAaAmQJsEUZbGu4SVyLlSVZFq5FlM
stv1pcX3FXKEfCT5Fwo6Ew2016XzzcMXzxDBxL6VoD2bKkXEjRw4hh4wVQAL/l/s4+gX3lVRpNRr
/PTd27BU8LX74/cQtjBDUaCm2Pc6no/5B1jhkdCwHBykvJjTvG0qTTu8dSc21nantD3/esDx0ged
zKBGuoWgjb34NOn2HPWTbn0DyKmq7aNwJL7ULAm1v86oYW3WHdRk/EhUR63YnUiNSgS5DHBVC5CR
oriI4JXYKjbQulv0TskDuXJMb9+lSlY1chSiyURLRW2HgtACf76Yeg+rKovbSMA0RnzexJwNQdBi
kwrtFoTttOsE5F0RSvrkJUh61+rmgx9p+VztlnZ+TVCqiACeFVwvJj5lH7qBnWjKDT7JCc0VRWwB
ijomQIOdUboq52FqP+/WmArGu6BFwFz5KQHjHASr5jKw0rtL7o1Qs93M3a0MTJsH6CzM3n/4s6Ag
9sy7JTN1d0t+4D12pP6Irtf9qpOVboR5XBHwShDQEUWD6iYlldwi0rEkKmL6CHwOpVt5MD3UVJUr
0Os5JGnA2CQrqIhFnTVKHj/xp3sPu4EdTbX6VGGv8fsYH9K5TeSFBlY2axirdKnE6vr39eHxGcpK
c/JJu9cqNO/k+p4vwFhovNK21AGd2IbtWBIuAESJAHrj2OouyVxvK8I5EXMHNcDgyu6HaSd1hfwh
Bn96ATSXJCx01uhuQRv+C3e7a+PRyuneeczVovZj5ozjvKm5WsxByzXfiBau0Tj/WTXOYKRu3VF6
wR0SNMcpVlOkh09Nd0mWqoU8Y4Olmx48O/diHDS69OcJ74pL4cciOUcYV0/upZT/fDhIiR8fejgv
bzTzxxYNJw+HQvMrsZ7sNvZtZiyO9UZWh56hs6tLlBXF8oyF4V2+vAGAhxMA0DjwlQy0pbSA9b5F
tl0WtYaHUfHwfRfvoq4Ut4IJHGAIWQMxwanSMy5lBpjcDLqzGru4AqVBZB/hUVa8DdMtc7f1ufzc
fKv7JrFvBNCs8synWB8SoSTAJmZ8PHr+JriVzresUZJmTADLHfmHVdcicfE7QdEo+5lcSZ4CUkdT
7XAj8c4XhX4N/o8phcRg6beFWBrl/0GqgqeL9XrZsRd2p6M6dAZ/ZIIXh3U2mpu67GLiqgQ6EP5n
TmCmPBwu2KnbV9iAAlWDQuCVbeZ0lnKhM0vWZ3soGyT7mdRgTdNGXqLuIK4SrpfCd25Fyr/5d8CV
/ksILH/6OLajbqtYmVuklfAJ2H1zm9F4tZgAm6ojS4XgHGFTvYT48mkQ5DdzD0LpjgHGjtpKoFM7
0roOml1xE/dgW6+/v3kydIyoXpCEDKK5F0hUB5iVb4CG0e+2oIv76QYGQJZQLTnX2bQ3SwkFKxzp
JbJSLrDIq2ULLGyqBMvN5I+3egS/QZcoF5sKUlUt/LE1qmltjdoiUodbGbt4Mm5aomsWNVfPQigJ
jZncpySSWnGrMWaodIikw+L7x8JgEapR7uwGe5dG8Hy3y6pz+5yG5c4LfUCyfeSf2Wn9Q9QVkrsN
9nnuPShafkzvEkc42weos23MY8ILcvySmCfs3bewAvKglCOWdrGPyWM7H9CwgIewPCEybgmG+ZoO
JRgh4uOzWjr6sANgeoP7Nx1s0P0k3S5ewfiite17U7WlHpXqc9tE5EN+DEvcv6CCLPKtVsDpLu/Q
Tmk48QQrsXwXOXG0vQVr9wY1713fud+a8gwvtPUKowqlHEVrDKtb1uz5GYcvxVP0LJSlxEQghVPN
1LG0pn2C3dDxSGDx/+7pi9yFg4UIfiQ5wuYV2ADvcQkAYYIEGNRL7WN7AAXNV4MLT5S+siHWq7EN
21roDP3rosKx6At5fCeqk8Y0tNaS7/zXEILtzH5yPHtW+EAoSVKRC1WuDXcLwwqOei2jOf8YsGUJ
QG3Y+jrJUyIYkNrMU1f5dtEHWgLe7Erxak/GermCZP05HIdhwHwNn3Dbt1KhTskqGqbpfbi1pzrV
U+b+VrRFcM5Mmb43hAttHYRba8XsYf8b0sXCagDloILeWf1fzaC1b5rxBGcTta9yP4bE5yXyg5vY
I0JDfDJJ7k7tFJawW8qEPGUwj+6e+q5wvzRsFNMH2qX5gxatVgeeJlDZcflh13Q1RlgFiHUYgER1
BO+rO91glGRWq/MIJjYEqgcXOiSdMUlaNB+/PNr/F+7UrruV2ZAsYEHT/zpFfHJV9ZByL2zsBrhO
nzH3kzUBn2xxwm9QUBSK5BPMWmae05eoRXi5uZJF5xndRs9EN1bynoj3K3yTS1cwa+mLj9jElscM
/iS4rCNr2lwlHZMmCVj8KvRDiuFBSJwHTzH0/gU7e8PCUM2prdjJS1fcL7bjVX+7U9f1+bEVJ8an
twSP1pmGdq8wUBhzYoIAQN27TIH4dZWVy0UT51GMZrJFureC3Mzeh4WxHTTHl5fq782AjihMul6a
m1AX5SqgTzQXwzmFiMdHb/D8AvLbXasuhalT9qYBhmT0SClHYinBM0xGLPGl7usIBpy18u5OBXpX
s76c+tFtUY01QgFakzoCjMcMOB3qRa6rfxc6QUUo6SP0VmXbB5LRqOb9RMPNE79jQU0FP/ILgk0P
JdFj5IwKaFRHfJXgwKwBeLHjjjwWvo/ceLjefcmhvMZ3yCq+wu19w2bkBOvgICmHQweYjtLUJGRp
xnmHbmteUGBTfXb+pAx/GssewLufG4g8kQgkja8msPXBUYwF4GZk7UBEdzKvONjhqxcILlnCDC3L
BAya4RRRnSWzeC2xgeI2vI7B+m8Ft221oGQhwfNt4bd+gq5/qWwMG/vaDmGLO+n/Yei9irp7BYDN
xgSqUcV3GaqV8uJu2i6q2+Nnj1wkan2rtJt4KOevAtKRtSZ3UyOTZCJ1RWIfQNB3v/7n7FfX1y28
c5Uvooi2MtGKDHK17wd20ZdtYVIUJnrFTg1jbImE7LqbNawkH3uZN6KJYNcweaiWIpVKpR4LW6oc
ouFburvyefiPz58xMRk3m6YGEiReLNrSAg7K9CmU/4ea4amu3kpjxUr16YU/XRkbNxYNSp0VD3Au
97Lw3XGZ1KvXcQACodNpKIefnxcO580iCZ/tj73GXoN3DAZMuc70MjEMLZCusr0dNxvuznKOtXge
gEGr2kQxJrdFR1XUUdv7je98D8A70trJ2zZMezGh1tAIVxiIfFxbVZgFg9OqtxOf0g7iVTv4p/2h
/PuhPbTZ03nocJgDeOk1ECP/2R97p3UGcDoNvCTtG/YR0Dh0brHWqU0C3V7X3l/51w3Z5yYXGyD4
07FcH7dnJaTExQCPWZJF2kjWgGB1RQYfP3dN8l1dYGkYQ5IF/p2LkeBw9XbVpcxSGAbGARmlrdZg
B7SIyCDb1gtHILlWgW6yYQR3f22sTD7KcabYN5bdY7N2VtvQ7k9JRczXGo9g7J2LAAc/f4TOMMjw
ru9dI7YzOiCk1aK6Oj2Jr3LlZ6vRez92Aw5V2tBRXFb4NPSdF/0fixp0v9KMCusTAQLR14ZoQTRg
hlSbfucTbC7coQk45Z2eldRNDjDLKJiEtWXTCHxS6RjAcyG8vH3wSvBtHm4E+PC6NBjA/7ssSWvH
PYHrLiVEHFQWgAmf6/i1nFg9NRl8ZZ4ySsuX9mVQwSSlpk6hwJAuDj8Ikcz9HhO49hlWI6CvLWw+
ieeR0kp0EfxYIEMWdVC9ilZ8e7rewuUsz+/eaP/ATFZOCI5D/iLCATVTmIG3wU/s9FDzCNTTn0rJ
Vd4tK5jQ01WdFxOI5AJtuWPAPOuhJwHapWilWO4xRSvUp3iBPwS0+4+e4FRyocSu+ricUVxEYWbs
esh97MhD50ys4rithiIgTLDUml1+I0hKsyoZH7uHjZ1PIxu0bxh1YKQ6eKwiMDXGoAdgoTb6KMzq
RRCiKgeoats0ckjI4zBJsfKbjajGoM9AsfU21h1k6GIoCE9I3nHW6ycZKXj5HWGpRaGvQA6q376l
dLQgtewzSgmY7Npybd5lNChp9/aOMglWP8R9Ue0HG7Vm8Q98Vp4dPLY+WLWEjR2Dc1keyy0HFtTB
02fp+oqxNyoL3D7I+QZYzpYAVbZ9kDZ9aA21eCwAMqwmiusLuQRzRgQCOkgDgxXzWZ3KDM5c7YyY
hRY3pDh2StvAtozucCUPKC94PohTlP0v426s46TL+5U8B8pcBmbFQ4/iUY3zrvDtXtGxGuZdPetA
YGe3InJiq3gKH5nxA6Ro2vgqEi9uyt5GvEzS2HO36pI7Qgy/r++do4Mg0+maMM5tnzxocQrgtaRZ
cAjKKGdMvq5p18VWu1njqXiLv/8+FwxHH3l10hiiRXKIKGfZG9lt06NMaYWxKkvqb9Tk10g/Q7vr
340EKMw1kMEUAK2JJ7fe6bkfxHd+6T6Dd8ZE8vghAE1FU8tYM/2Fz16G4uPAU3WDxKmM6ye6z8+4
T6w7s5KFHfaGZHL0fAJrNlrWLoFa0+1HWymJLCsr/q9tP340p+YxSSDMIebWtlXuEVDni2/GUBND
yoAoK0xZMjWkxq6XRJTh9POpme3L9a+XY4jPejjzAJGhyIBCOypg6VWZjTdjJLubcbZb4A19fad6
h6xc9xh3VYDEgFozT2mZtndyDPJ8X0iJy/00zKrC5MfY9EQVI1ZtTaMjksGw397qt7FqMeG5YujA
3KKyPFM2E5tlMrUYYcUwflUlkuHeT1R8VhV7VD4Kal2uymrFzX4a1ud+MkK3JT1sO6YTfrYmBI8E
gZ9cShGN5WKMpAM3uUvUENRyjGAUhRWPoEuNFmXZoCPKbxev4EuT6BGnM2lA3rJHWFGbapzG/R+D
7QsMGfGxSjkZFII5mTTPlIOh1gDE5hlbcWlu3cyFC3rgNx/sq7wDfqJnt1NH1Vn2HQQQM+p117vw
lwTeyj31H0A9AHj+HMGGbS82kx5ta2J+NNAqTQp1MXPwMkl6Pl1ZIvClsPMkUHw3qJNBFH/hHk8q
MmyvbmjHHi5DHx6E++XiBlxBu+m6qd2BNrerKSiA7VEMaSu5VGFye5ehNa9hKGzQyRBNcflgFzKs
IJK5kt1a1O8VR16zmW5+yyR+f+FkzMYix/CeCcaSprzPcQUUxKUG6/LmJGuKeNzPZf4D/CJ7Uh+k
J7KTQk3iB2DPgC3B2Trfh3fpx/xT8CZ3QWXB8XW2xkXdDvyEEO36HAuzmq+fOaOw39ALnyJlTOJr
OMB1SYhzewZj5yzWSq9GyVXAKMaq16vzFCZ6cxVbqiykyqObRHzqt7DZsZeNnJ3mO28TTilQh94V
pRkyhX6sX0L5Scq5aJPlwJGDcyO0NPnaGdZQyuGlVy386F4kJ+DL0ijgz3k5M8kJw1D6z1sWt+nb
zmi2UAwad0uwJAk9nw2+7yHSdBQSXTykyIiw/uOtoCPWMy9UnZA/E/FVnG6T6uMEqZ/7YswcKpZ2
XhGPKHvPi+G/xW8unUp4xgGT8AiSqvqk0IgaLD0j2F2GSaHOvTdfU9hHPy4hnm1omFao8cB4hiuu
9NGCeBUpTg/+0xf2Pk2C3L9yyNqTqup/bHhuQHqFDxsxhLGHkBhw/yf2fltfKTE8x59ZxQtxElyn
CCL0ZnxaT1jmPsCiPfLpWc3penkVtLhOJ/TAz+ZY3K/P8Zh4KYpCch6nn2QKipAKCfpKBAGT03fm
ObuWK4fdHBsnWvtUd06GmGXhHRtKmqU1JvjPcK2AyqVDErE7d9GDEydY2YhQx1zLV8KFfyWOu1Ln
R4/SlUjbrvUqWs0gWSbdNOmNQgjRnNICLiwR+ocHVFd3oVQmBRUWYAvL7NZmSpg/mVsdY50aMWdy
epXVwHYL3nj6mgCT/n0bRa5xjCvu5J+viOCQ4DKK+NWlBEX4SGV7r4UfGcotZZM6eSZjPko54qTf
rEyWa2MDHwa7la0mK3yMKUKqhNHeqhvEvzzKfmstFdrK5GMJrX6sdV2iWhrkwCuERlyh1OdkOKdo
oLHAy9ZS4J1gcx/7nY+ZbmNvPL8fAqEJJ038nfdtHhucTNcyMfLPD4PRTJxbxFOjIZUPRrYwk57y
6lpAZLPaO0tRAt/ZMnyy1Egq642FlFUpd8ahZFrQOMPbBbXfE/kgV3xstQw7IYeYmsbZPxDQoFaP
e6ChXsFWwrTKQwpziGCswemjWubYeVYJZuESDnYh9tgm49hfhg9jbg0zRQdXsO3KvFb8jVgHa5AB
oPU9+E9xZn/Jcifg7Z+y9o04HgsGZCuxrq0FMPP3kmvxK0UsUv0rIFgch4faqwHy1+e4co6iSzfk
/ZHOaoja7NukaMTw35KUgI5WIZ3TzwYYA+wIafqeUZSlrIWpbpleOFODd6BbIUqGnuMGXtI5CCPE
H8W2X+Ej3BtLo4iiM4GrlqJr2ZfrBtD1dplyORyqgL4BzCBEOSVzLL9gJf5/4kaC8/o1hFU5okjo
rtMILfZ/hyo+2cFXF8GOGzRLig9PB7CKhQJMHZVmZDAyQ/J5VZvpB8f8h1TQeJsy3JIaB5YoTiaG
1OQNMZFpiwr5m7kWfZCHDbyvLFKQIFmVpOvdr643KlsWtOWbuwdaGOODmUIvXqRTCBqBH3HWCLNK
O3JUKkBRpoc55rWBmXmOQhAlpmhPShrNLl/FtC8nyVZorMEjQ236z/gg9eJcrRLzEFAsaM+OvTIv
i5sK0YVaEDJGhtotoy1ZWlPHTEO2lxFQeIy/wW3HzWxSw3h/qnTFwzua4aNcuZeJZhYMsMh/ykhd
ykccJOGtc/7F5b346/qC5pe2JqWrD4DWyb/cHOWr9jtq7/8MNu7ch7TjDbwpOaP0F9f8Iygf0Ebo
0UbHWnQ/z04yIxCyXobSMHTM7hAALgJ3nooaEL4jClcvdydN4HFo/kd/B5jY9BnxQGYPl0Zwd+6M
RT/LEZ1qWCLKXed06gPdGLMrOjIBorMnQHfaUPzm97+Gp4/ty5rm8wOCuy/Bv0RiyrF9ZKoO9KJ4
haqdqXAaEPTbprDTeOBQx6FWKmrItv9aE3stKh+IAtCVNppjaq6SB7aHEcLMJUPNnO9Gtd3ACKQD
Gxg/4EPPy20rvSneKLiKTEA1rhmCTRadp+rtMtrn38npso0Q/Uv+z5TcIcqoGLCQGb1ih/rysSju
abW2MzFZ2lO0IMQr3MAMtODzmSuKxR7SEPBalRwVu3JZqwP/PfQgY2zI4DjufbZ2Um1SVeFXPPrJ
f/1iACsOxUQ6UKT0IlSraWA/W0ufRQkRRlkLcxCc1AmIuZtxBLITsQA1VCIpsSqphkHmxx23FgE4
gk2oqZ+Zov/IFYu0VypIQXyRI3jbAMSw2bMrnSSBWSJtcEWK6R9/11FwTtEpsLuSHcce1xtofCpb
iD0qtt0plkB86yTQ+YUdhhNOO1rr5nqHGkc4ZU6ISvhvY+Igojy2+7KsCbeYRhK7FqVWsY/cuxDT
D+SWoMxt30MM1MlZ7ycpli5CNGCXoMJq+b2svA/cTVXRULFgWtWJUOWAhzwXBvquPKTzT+lRcAtm
5/6ZX97YjqXEAGIWMzBg0SSP4QYE4ZRDZwvOwaEztrR4Is2u1K3dKKO7xVAoffX8lChz5rITH1AF
hYOGcEaJ/U3FuclJsTqvC7tyxbyrObo8BYelFqppY6r0Z1vNA9CsLYJBsnS3kOcnL3hIWnpyRhsG
8ErOSxEwclfUhdeJhLJt33LMQQz1OcT9h2Z3t/lRgBOXVEWkrhSkBAp/53WZfdtL8u3dK07FMFe+
aLBG7vKIxc4l7VqlFb8D1lluUkBCKASDy9Lf9olsP1yKhbjH/MseLG/RixhUB2YVnlvMPUbYKhgT
Hk/STyU5cFwoaQsui/2u2vO4Risw/joDpdfAd0IDoZN8jU74qqykjPk+JWuDVJXfWiVwgLXszxzP
LdNa9rSoEH14pvnpPK/OSGG8BPCtKjE6GjdmQOd9iL3htMaIxM43llXn2yxpAcdy1DVnWZZcF5Uq
owz5Y2aEox4zIJ6sZubIh5FT8CeYOBviaaZu5Qzj+JLVJ14SZDjesdprGT39A8Bhnj12x4TbFmf9
2VCJoKmlAfGCO9zU5s31Vy5myTbbVdFXBNVCbIlZ6rewf+59v76IsMGEAQnSbk5Rd2QeyNWt5bf5
VDDooKaDYpnAwi6LFTGy+vC3oKXSXRISLqu21mGJRGnBYrCFPLUB11To76UUAeNrOTfojT1uQ7pU
J2nxqGrVnu9zOhqJV3yo4lcbcyrt3nsN6BauTEIjqeUtLP4niZ89Wwu9ZKT2JD9i+3okwJ0HLypC
YbxK/1+3+Bo4OlLq54x0T2PsvzTiHmwAaJgk38pWe4ivfOdv6hmR+7oIOWMBYEo8vFXfiifQY2Pj
21V2hiwOthUQw/5viXzNPk8ZuQqIcTvjQ3WpnXPOIF+3XoTREqbp8Xg8S21VGFERaRg44EVt8HRW
FZH5y9twMKwoFDpbCaNdXjbsSCKP/ixisK46IeDCueVSVXD1l2FMbMbIOhCvG/Xhp8OxBSEn5bZj
8x7WLvnUq3oCnMNQ6hZU67/SIx8t7E4250ST8oPyY0G+JVFZrbuU2KBFhWwxLIyuOKFIqbFGHuTF
wDfVakjvwCqbGMlqw0/mOsBqkyUI0tjwqrrLiPpyUiLKhiCArOmI9wrZOoiGbQwThOMU0mz+qQ5O
5AygV/MMGACWSYqX3cnUcoviujanGK+LTfpkOlsvv+L++6Yu0IsjQhZsWK+Hw+Tom6EtWm3QNeQ1
zhUGgtont7AJjdyGWu5GaqhN2zVCSCWEZ9uy0pEa+i9HCoRFPeNYrQr3fS7omu1Rjp+RgN1il9tZ
zLGrvi2t2UxEOT9WuO+UA9cVsbe1jtli6D9SwX3/3PZuWVYSUjQo9BZVuG2kSJlMRb1SqsRcJxhx
hHhkQP3rOo+ZhJNVhaHAHMViEfeTy3sOZD6R6z0H02VwRxCFx4qCSsuSX/CceP+zyhOw1Se3f+6F
ytwZNK0GmnBHxMzbNu0RGuR8AzUeTM1zBd+hPI5Yc7os8sXN/ojw8zK9M26CGAEuXi9eybgxEsuu
5+DYvGZsAjEuEF+CsWPodBt0PJx2waMOkozOcvzluNxemamoy2ThghEPHw+qknlqrCcjvV/Wk+XQ
qRnhdfptrKjtlJ4OJsv+NMxUMqVyo1xhyJjjGig4/XxZGC6zTr8mmA4725hc+SWGTuZ8ZgKZTuFW
bUmLj2/JXdZdtdgIC69O0AgUO4naXtTb9whVWWNsYjvkYP1TY6mv5j3rDIVmwdrR0cY8zw3aDmXI
BvPzJ4Dh5QvPhLrXVKO7N1njBnOZaxCZUxbKZ9oSCZ5oQb28Z7IIoWsWVSxVPE2J7aQgidHOEyPn
XAjK+LoTCQmVx9O687L/1FQnvZ9dKP/ko1HrbIR53BNGrdK/GsrkVj0KNkGD8rBTphDVK1nhBWm6
SGdxplaO247/iXJs+f5lDZKL0vRLlniV4zP0SblTSKsn4SDNd3ZRxqOdHzZHHZgH7QhobDbxVoF9
BR8gCeOdWm918ODOZQH9AKRjB2gnRfOmZjV+eest/roH096oBhyQAqqKYBb7+iQ7qMAU0lEKIjMb
RTnVa/4iGlE4oqo+8r+N+aDqaK1Ezvhtq7DB/ZYoLwZXeXJ8Wucgqw8v/ILKBT52EkFX1tIU24do
a3dpFpfkxbCIi+lLsjWbDEhCrUsEq9tnQ04O+wVMy0WUsWZiixJB+sLSywAOvnJhwstLlC5AGU1W
cZK33HMCbN0VlFsqb3a3/wKbdB6HPGkUNWjVVnQiEvEAqC6hfXQUc9BHx5/JuLijSzo2C3fkH7XT
1WUr8YiPRrjOclyxgIoMfGDHkTj00mKPSrdU90hj+KSuAzFRMj/hBYXSDyT3S0Dfwi4IrH/4DxC2
nlZqqF+Xxz9mHM1CdZ7/vbqQJ19RCOdE7Sb+kNDSA0qN+RQ9/2DHAWM1h8su+M14/brXhZ+Ux466
kq4KLV3KsAfgvQX6zE6aGa+1jB7Jv6eq9ZMOFR7p6SOtJoz92M4/QNzM5ewbSgkYKUfSqMjq4cnE
tm+ISrfv8AQD6SWxSw6urcXJ2eyTkn/ezgvpxHehwbI4sWrIKkkC9nluPvi+ohhuHKqwysNI2HmV
qNcLk+wUduczV9qYYRThulCs9op/9PbwX18Sw6lk9xx9KQMReee37A1VyinNc0yngThGatc5yR/j
6gg4MM/8vTQstYQzyP+fyBgjWTFSn4a7OgHxNqRM0Q6WDElcvQ98b9fXIQGIgHXTQAK9AohdA6WR
p2s6J1vsAH8Vz6oL0ov3fOlfpZwJ8AgKNexw8k63eVRNqwe88YrRfOjSYubVhAVay6wGp/flQHIy
kZBUFZP33VaQpGIgqMlcDHZ7AWzk4gywnGFvPkEj6K/z7onbj0ERvZX1WQlIvNemj+nSsqY1i52e
cQihSYV0o/OGYpOxSBRv1x3Af902diMxgfyvGo1D+ulTtZPcrx1pXrtwsl957CHLnWMFz2f3TZda
0zGH9ImmOj+cqO6ks2A5BIU3C4TBkZHlSuLdoBEJm/GHhN6BChX1g/q/KD2joUfmbjN6+3KdkvOA
3iV4rxUcFs4MnvJsIaC9iii+RgKSF0wYBDFvZg+YfxXkUM8B1ZDtb76lhz0ylmaLPjxWPt5uOt12
axu/8SgRXUhj8GfYZMGZdtgMSKLIYtho/e+Didgdfm1tlVfy0/Z+ZPfKpYjk7/Dlk9yx0oziixOm
Rj63NnAlKn3zlNMb40Uq07+yKgbx2+CgxoU3FbMu88SoRH4GHZeI6St1iti5PeKwPuTU9oeE8/y2
jEcogDnFBntGNh1LNj5Sxk3aQ+IAQ5boUzjnzb9XpKuSOcHglUx6P0ujPLCVjly4K1/ztXvWDtpF
o4VAzH2op78K24Y7RhGDwnbN0iJGSelBUfOY22k7lL1rQU1F7Xxe1Z5i9DBJgLPMflQOqSgy2koo
iU5FdAwjgC8OqWZh5fzJExYzLFXvo8OGyvPFspY9Dpr5/Czktv+aDwQOUu+s4Ga5zArsMyOgUZOZ
tj6eJ3/in++FMlzQlcSk2Bre6JwAjbAyt3qnftdtxO732Q6RQqXZkWYlcpTSYcWyte1J4fijKpHC
Zj7eVfa8p7EMe6idaWu8MEw3JgtFscOByYIdvvtSfooW3IKnqinq4aoXoQF/1ESdL/oItQmqjw82
u8Se/7CbQz0Qkqkti6Lf+O1vSpOdtlHO/y668bX2jor76heYrkTo43xGj/I6f8T+v7dTbmsFI/8P
t0Gf1Ia3SHQm3wNkTfzHJD7KB0zNeEj2Ywc6HvKglE7XaObs16jz8Ezrch03aKfrsctpEataUPF7
+1mYY7YM1vk4f1N1Wt3KLFcebNULeJ/+bSNPkNEErGQXBkyzRFwUzrTQUIm5Iyd4IVAF9cJn+8hN
qWXuTEmQfY1j0iv3cVhC9AqJ5OqGS8nAYU0rdX0zggjeVG9vOeejIOpyKR0g3KFkbHHR1HK1qldB
O8prb4O7FCXwW5fNQE0K4feCB6XYvqfdWLU1cT489DYrNTYVcFVPTIHE3v61h2J+IWlzbmHOr3yd
rB4Ear6XPQf+C4K9mT3g2hyn7G5U2vz2uDCX/9DSnsbKsYGeE3RRMOZkT0m6UAwyv78BpDFdkUjE
KTdGjwldl/lFZ/6MsvGQVdb6pJLvILopfzsXIUgg1GAwupiv+bIbaGu8rWQnpPQBDKtyMyzcByhv
Qz3AEwIu46534kEBYejBf3r/LCmcqFR1rVq+E4kBe+ug/i4B4NAq8Jrb96OHW0pCjlcSPtKCuFk4
0P4PtyB28BZKt1VFWk2am/ycsafgWLoecDNgONS1Clxh6RGdInuHT2WOkkerv67X/6nOUz+7kval
oW94S6XKp4dQ3brtKtDRG0fjkLObxABkqMvHAhQ2Ub6OZl1M2NAb3RUHJ+e+RjSyscKKXIocJs9L
5zbS2LeO+ZWyTZqyMg2muP4tiSODwGlPFAjKiRSqh2eE1X4UeevPiaKnX9UeRWJACLPBDNyAypI9
p6YfV2U2tgGwDJBOlHDQ3rir+ZOCI67oucU4omj9yFy3D3oQzEqkVY9HqRR7W1FuyVlccyS+PG4c
3rku0+eruhRLQNesiw8lZ0KfisNrCj1yfmlMRA8gWm0SBd7IaMOcvwF1UIgNi3JKDOx1j7UQZRRJ
3rErOTpmJInfuxaIqoS4cv5RURO5tYy88eSsk29Pckgg/A0BswjZx/c3m2EzXvRWcv+jjG1oHTBc
jXnQXkGdFQIY/ICVhFFgRIQPvZD5i9UWkpH4Vm23Xbwc41lbXKcmGlnopEmTL5kh9apMy7GPxgej
SqUq4VKP5Ne202quJfF2j2sfXNxUOpyiyQhvyuNcwr2J+6JnqEPPAfW/+K1uqrw+8Sdcfi5dsBYn
16O75m7VDlljXhwizuvJeG5pHBKhn1+WaXf8qsJmhItvwzQmAcPKhv29invpqMe5NXYdOREro2u+
Dr9+3U/8HU/7hFLvlX1zNnEaEIe2g7ZxGyWBb7UBy4yfUQjrNwavbJMSb25NnTNLmTKjg/5UuT5y
v+krx6c4reb/rLSmW23Ft59lKBEe2MreKWOstNaDotKVEIsMkHDWzzJDBsB5EzPkcywwAxYz0HJE
gowlueI4qsO/42PA7AKAyQICjAs/EPqDt7vKGo51/tW+jL2TaP0gFBPLS189MDLvfl0ApCKcX6ch
j5te/Gy4fU1zHovOlgdLKA9TqZsBuY0pWIT/S5/piGGM0ZioC2TF6/skVSgKW7bGsni4XDSXa5Ld
r0hdRdAfvkf4ISFjZ6e00w0tLTpLNeEdNo/YedhEn6AgmKnt+HKA47/h7/+U11c5+RscMKwHlilz
pKgFfpta8uNYXo2SyGnD+R1NyglQu9kkhCrKnkjvXnP1Rmm4YgJlUdTiXZUj7hTE/4rzfqgWroSs
TWFK8K1acPkVKxohMYVkfIgMNIczFoHHJzAxU377CqeAdr8gocA/Yk9R0Pj61H29b5OG0yKyaO8x
kLFqkb4TObnxxgSfIAWHdcyc72Llvqnq8N/QVHJcmt5uW7cOJZHd82yz66ip1xCrRRLdYt/Y09/m
TaD9u13Tu4xqrIeKr9XfPGvMHYJL5XEBH4qFEAj3FNC/SnSx44xmLgTIT9Z66cTniUozCqO2emzw
RLhSGhpw8wLz2B4DM/FtsdcZTaDk+AKUG0GwnOnkqA9jQFR9oViLH6TCnu/jG6rfLlQ51K2nfgnC
hYFovaYHIADcTuw7StjtCCPngbxyB7LBxffb8lFfAyvR/Yax35Qb8YwVI+OBFrmFKT+NLcBaEnR8
PcRzLz7c+e/V6oOzDdWPa0NP67tqP9lp+GLjw1g2CTU/SeZngt1uULjaY5HO36f3g5kRyXXw/y7X
SChL48gxKydeOb73Rrafoa4J3aN6yDIIyj2BzA1o+uVy6lK3peDvvP0jhibENfb284IzFa6cwx6e
+bsJ7aB8wp4eZPwaPCfxa5halKfTF1ak4zj1uV6ES/udxTz3X+E13tjRUSSwUgBN4uk7PYZH4rQ6
Fpcl9BkDaBnA6AAeBR8cDXI7bL/OiSUhJNdgynjYFzc2QeicnNKWLvsU6HebxsxwDST9IvpFkni0
+qQuCzUav9F2TKbDX2nmBKjBIMvuOh4ODctgBlcvKWtXn06UD3FWd0lkxo2dk7RKwJMS1Z5uGbYt
Scx8fEOVrdG720uxTAdFf74hbD+MconXqR+Fz7zaZ6HSXYCsTK5NisqcUjki3vpWYq84kObNJy8r
p2ecHmyugAmWVcin4nGlllfNoYBWci/yUFN3v3QH6J9b2FsBwyFDx2zAC7UHrBpvYgewevoUghAa
QiFCow+xR2JVWGS0O5a3d1xU2zvMPwkGp6847oIYsWBG3cbIslSLagcaouSJfGI951KWxIsBLtmQ
ffYDKuLkF/qC7AXiWCJX2e4guzKft2M0BzJvQpKtUifru3jUO+qS4UWN+tpn6W0QyDbaMMgz3mgF
pgYvLEIt7ktwac0VKcbl8Cz3xRi0lUomZqStg3Z3qk9eeoG9w4pDT51ycHctyYOOrQrw/N2hK664
xsZXJhWOUPUEVpZ0qB77LQjnNpfD+RYOGhJxDCvNRC8oWQbhqP5bp9uapGPYPBn9putNuj/ubrf2
lpnpkm/bSdXVhYJI6uivP4xqrLDh4wXaG04IFIUEDij+uZ7zrwRHIX+hTZbkPYduSx8PWtBktc3o
K56AjOXpAzqf5Eleg8ymHunIx5RZcVkvR4poi5cQX+5R1OogVU+aG4iE6ONqDX4MHAHpWkAUlTNe
HvGnaXl+h7G3OHFBnzNaOa3JQdwbs+L7UfAtNtOIN2kIg541KpfZ+bB9TDdTcZWvjcnGzyIFtV5W
VrkAarsths75M2+BKIevj0IFQGwpqIe1LMiQQp/PS+4mdMpQsYASqXW6wNzGSwtRogMEBEPTi7Ta
HXTGvJziy8NQ0X5gpzA578U9sCcRKpDXRPPFOOX+P1Fs3PbxXXScKiJOEjZZDmrvW0w1XYQ2dQlR
6e4wPTMJmKXQ0ajzo/2SZhpS5p6YD+81vSe3CCfAeQsxjbWJ9aigLlZjtSTkLGFr3K5lrBB0x3ll
MQ5HgpUZxShPPFmWT1bzhDbt7QBzIA2LlQa+vkLN40Rbs2KuVYesqwCfpj+2G/7wB8YQF9ozoPWu
9QttHkUFkJiSYrG2r7WyQwygvUMN7qMlaofx5CITwLijG489CHVys3AO0+IBVorYp2/CF/JIky/e
E7+F+oMxswD6G9DZ3CJYAfZs2UCnHJSMXFF0ET/R7xadzPWHntQ0xhI1WHc0U+WLoY6P4+pYRgaO
1HhbZYaxk4OF43Z+fCjLubfouy+3hFK3+I9GE4z6YdHOaWUFCU5S3DiPekrRAIlz3KQ91tYQ5EZQ
tK6a2luO+IpxMaAmLMWBUl2L7iSijY0eQQbt64Nd4VnlXH67kZs6c6Km3vR6fwzWrISD1giSU2Oo
zZmp/mxvg3+CEyC7FjAHHsMvDSN20ifDnxhSRKXhjAOF+mVCsxrtiIkGBnbcQmmfvKvHW9dqUBpN
cQM36F/rug8dr7H5/iXPTd6GGuyLBr2CtgHy9CCz/oR/4wUpGw54Fj3R4DHy/kwetY4Ed4UHYmeV
YoBIDLnrHVquYUQyjBrhjSU/AQspypAw5iK40rUh5UNItRFFFi0td4SFV0o0w6eouHKiniEyEveN
yoO/He9oL61aHwh6N2f/Iq+qpRNnla0ZfhsqcSiSK9XZsr+JElZ8uirHIKj+KKpRzwFfkqumb0Nt
3n1JfhEPWuCm1JlK4nsQbzmAVXGLahEdbAK6mkdfmTIhBTwl6Bi/Hm8wITAq0FJwX3E0Pk9sZWbx
eylWHnu3SIiIW2awOARWk0MwdxqMkbQh6CHjgpblti83F1DS4tDnjrSEMIOkuRTpKlU+6ndy91AX
xRHubxiKX+41tt6zrE/mN667gks/A2skobZb9BduyFmp1cE4HrAFuhGEg39wDpayv1gHFkOgqo+i
HE29EoWuZ6ErQsntQ5W7GX6CVeAqNBRI36CCOB2A+zqrWpBMPFJLD4MBoXQpe68FnWgpV5utTn0o
/FVKkEqCz1M/BIzOYDTq/6jtRyTLz8eE5fsaa6WAupesVU8kiQrdWpjduKB8gAG/thwbTcFQaZ2O
ziHLBBJ3IUChWRXADJSWlc9Ftwgz0gUzUXdMWeP2wB/gKK13CkUk8P951A0OY2OWQ36H2J86098G
kdkkmDE4maSIJmZg6OGu0I4jDpHxH0HA7arHlhE7RzMnkufZywYRF3fPLhZ15+Ty07f1BfHStr12
RWtvWSOOeBM9qCPx8xOzSvqekscNbnCh9GAQjdIrQ3FnjI2St4NZGzYF2/+W6diF5POyzc771+WL
Z+2w/K8DuqLb78C9vEplV4KsxXQypTJzTjMhuYxXVVdWq2oqYA8Gc9pPxZFhTkOuO4B1RHqL+ksY
FF34sXo+lTJhLO6ra2Lqd4c3NqHoTUI5ZPUm6dQZ8Jme8ChPtDb2VU/9kLp1CbZWZIQ4KU9dCdwa
OATk1aTi3na4btc0TtUCt4uFL85DiqvPVAHWabEzUeP0n4k5E9rPw2Wvg0oN0VqrWtV9R0V3izfs
MiyHp+wLfsn6kjagzcNGqSj1aMbiFVpTlXYkoQDrc31b4QDbXzQ/HY8Gp1lJ9bgYlAsug+cSOk3k
YSnhY1BGVOFJyp4e1AMg9hzHKonU19C3KhAicLG/lB6IFyeQpVL5bCj3Hl2x252tK8wBuVeeZNM+
YIa8xlkDm1iuD72eAOrdNLxcU+P19eCSBN/1aXC7Sr6ZERO/b61GGx2ER3JEtdL04+HtVOki8nEV
hUJa/6KJgxE6k1nonZonuKSzGuD5t+VMBsiF4eZVu61eAyp28BDiWMG3ZhblQmAlEuBvoWMqS0xx
Mk4tKC7Sdb6t6BFV1POF2eX07fU+AXe0vH/LptP8JFcNGupZ628QJ24jtCce6RE2NPAci2D1pEQ0
xWFwis8hj7pznvGlLv3lLOLVbeG6SAACMOrAMBDuEmhuQVmFqtC4TGL2681VpUrQzL4z7pWPFC4Z
LT22bAxBNZ3/geb49dQ7PQfbq/slUDSaLjfem1rDiaGu0SNAlq17kGYZ1aZ2NTOQgwwc5XiEKCQw
U0W4EPcJ2Aw5PY6OpNstXRUDoNyFAkw2Xj4kxyqIi+dIptaeNamJ+jDnP0j7bvWF55lRD0ky0FaH
uEMY9gRgLP2QxddCoUjA4wZuGtktEyyx8xuGnttBYh7V+6P4eCedb6vzqyrPYxuIvaDRDas8Jsd1
BW3p8XkoOcXP7+/fhJqc5qovyHv6dqVheQeDbfJV7KaLdAuwflfWBLehaVgUB81whrCzhMEvxzPZ
s9wfnVTQ3IbwCun/uznNjIAogT5LRrKRR0798p7GyvdxA8Hvv6rU/+4le0/nDcCAbfaf6OFbhqXT
UsN6gxiqKoJaRjntHfabcSD/3Dba0+kuk1wSidqqt7aYeDENoQxXiCQmcjb+jA6hGyKXQWihzPrp
cmvKYJvuKafghjnQ0IyoA3A+ezI7EZfLMh5gvsNd1wEropo6Zt/4WMxg9X8+v/MKDIWtZksSjr8R
0LseBKsScjQfmPrbwvy9q9NT/oV8y/pDPhwDSfyd8YTtgI+ylOQ6qat5KK+AOFqVADplm94vnr2d
a+v8mpADroCa/kGqOnyOxyh1ccUivdDOkyYOGBHr+QHP+73x3ol3MtGlkjcraxxYg+AFUFh1Yxjl
mAn+rAFPV46gn3Wr733WQcF8YK7zEApax+jp6QSvJROLzB27yqDe/yZmSJ+WuFlD5HU3Z5Wv/f5g
UwcjbTrMQKjCnKqPJjl51iZzbZhvoWUsvsJZbE9QBzpPeJeps2TSPGQiIqP1hfAJIBUNNcHBVdJM
f+tOt4Ddr+1BFWXCCss63P+fuIFaDQ706cN71qbGsiNAk3x3ApRlSIvx5sRrEswYj6IzOHIl5zEX
1BTxKNlubkrMvOJux8OXm9Kuh4XDT1fW9kmle1WuVfzURvEZIeIzm5jBTcE+LTbxpwFyfAd4fUD+
nMCC6yJr+byYbQSGVreDW702CTYnUQ2Fj8wg8ItIru6c09TCZjs9HrLCcNWVmTVMJqlcRHcA3rYJ
ChQCsr/vIphZxFzLCmoUOzKCyBnyak7md6UpCPo4FJdQJZb1BvJtzjr29aTbUUQJvuVbHQsIZGL4
d7euMGJC/JcyX77bRZmVvqwJLDZtBlek30HI9ogSDthKUdCehgtOyD9kpwGQd3Il2+eCx5REqcHp
BlyxHh2FpxnVW/4ZKSiD+ul1CnXfn8JhFs/mWEpN3pkapBQqqcJLpGAAfOlwHXN3z8SkTHoqiYS4
+3kEME60eVjtCo3y1LEw4dJv/VfsCkDMH+LgALkPQE3vDDdnVpByz/15R53xUfUxysurQyP4s2YT
mT2Z8tQ783qmaPGBl6R9Vkskc9cBAqJ+4dpxL+U01efEGDRtmLVlpKpu+YY1l58sf77/tPtdCV70
Or8ZmJxwHXD1yTfwbt5fjm+5Gg/XT22/TsWHfnc9xhpRPyF8t17N1FJFUVtlezh05slVM+U+SycS
MK3e/siSI1KTKEUzrLJko51qZIxdECAHZZMyqcR4pt0YFbdpuVNGG/kJiEugKKve1NUuVKkMn6+E
3ec9gsjtOTHVmJIzIDvWgXop4WICpJrTWFzwQW/6cqwK+b5scGSur1cZBjBT03oohG/Du3TuWRZy
FQjMF9YJCZqzozPSEJWnKFMxAZs1HktqHYdQBNnijo36hUHp7ucSpxKPh9cv3+r+YJtKHl9QNKi6
SLBSuJPfiNJX9DRc6eOxCW/BBBt4QtcPZ3BtBXrXQ7l6b9v9FxdnZy4eHfY1f7Sb4hJUzOxpJDRh
cqsvp0JteoV0BxrNR2qQyTEGPeAHCkHIfdkK/VyFo8dseN/Gzmh85+zRaMos0rjMUw7X8keuafiN
NLLjDh/z1phggavVTgt6ZFqDvqTI4VeZj0Ko2mbr/vP2SqyMONydttGA3wzliReBN9fxvS2lR2ez
LlYIqdkQQMFNHcBWcuecPvPJgBcS7tdWvLMEL9uMt/oeS6zZ2DFggU1Oz04+YRyo1Waky+hAbJ3E
ZBVvKMG2oGnbGj+3Wwdz3wSyEDBEtePTISkHFXFuU2EJEOrEyiK9GIwVvFhALoE89rjkHerRttsI
0WroELi1osvTLWLe3gI7PVm+dzD1FX6hRY8H3mtenbPKVbeEoB6ScdviihzfFY3ALo1erPJw1Eii
qirq6ngGR2QrLIWBiW9Guo9IaSx4oXpk43dyNWH0u3//fs5BNaIrwRS0KTNrT9tc0NTd/P4hgpi9
pNwtgU0T0ider6JaHoRPo/LliGmnCHSlsGQ65wNxAwr/z4tsFhqm77Fkv7uo6Rwd1kqGrUVKmpPN
pXJ+H5h2FiMebTg9RH11lZre5UWBYz+3N4TBAj4mwsGY1aVwoyoLzEAHhYjLOkV0Pauk/o4BZwVL
ihnW9yguPMks6eRQ3IHE6JcyXONdV1VyRtY+n6Q6jvzmXcQc4NzdTIQ69UlmJmu6WAB7sdYyEtCu
nBLOZEynkH63ANz9ztyvx80Ec7qd0r36eoU748nI6l8BGAXvJcVVx0i/DT+uSO0lKzfkCZZvxARg
ARPddCaEwD3E0ooWCpE6W9bdBQt+cuOzk097Sd2wWyjXXEUMETnWOqCibHjglqb1ZlUhASXtoWzP
4PvFmjqoipmcpr9UB+gwy4VyJMZK3xzzsJjUNXi/n/l3bVVJ480qjzTpCFZT+F70/a5KCsSYi7vm
ldMB1L5a65hzmoL08kZeVkr44rSO47pOzxmxjRX1t7XCQOlz5AfmihnVRubQXvL/CnUx+tDVQkGr
P3P+02BmPIrrxPI/B54Y5QyMt+BKIpOkrZ+GIfsPrCu3cJTKYRooazxUtodC42f6Ys01GOJV6GZ2
1Y3G2/4+aVD7cnYAdhireJ8j1Q9gEr5kE+JySZssTz4Rq7jAnXWltxz2oOFgkjn3V7OGtFgznWX/
oh9WSenLjJtmY69kPKPrfiXCGSIE40EtCCeUSDEv1yQU2eUqxZoiUwab9bETO1ah/l/2qd5HKqI4
eXbabsl9XcdIH15BFoPg7GXR2Gt1LF91qUzgIsSTCQ2tRtXKhVJeZVAp/hwtqu2Mq3oyJyraeXnw
YKTZPrPYUDi4bcmDkSp/F4YFdGU5SF/wL5yH3kqO5c6I+d/SIvPr67+9hfLneOP+V9pvTt7H512p
AV1JCtPBot1VfaTM7gASumN4DDi0VuJHbfbrYAVwTG7+mPQXFp1FkIhApQvbuDCWnlZ80a+1iJW5
YGAAHLUTQiU5sDXzM+KyicJfd2eWudmaE9k5qEBotvYNHZqmNR1QL9o4Yg2sBrMARk7+OCI3yIUz
0bHki2IooVQavYH9Wji6PrIFyUG7KFLCAW07294t9ZInbAbrRSfn7+Z7i05U31xdpAFbE0iKXai4
S5fjEUiSLKcE/RyhYbJNVy2YuJdUIXtAK3vymoujahWcRrhwo0ckae0EYl2SzZuPR1e1oQWEoaKF
byJaXzY0ox4jLeu6IoxO4M7k5PrsgWkc336zukggTi01OknYwQ6IY5qCiquOgyQ6Fo31kJMjR7Sl
z1M8+b4uZT1Xjz0VKVuCIyT7QHOvLGIHUlnBswAIgLTzp/PR+X9aS2h+sr+hpU3+rn0myYwDLWmq
IfnfJZRYUtG/U9pCyFtljKpxUk10i0BNyiVl71TIzmxXkOUExu4SPPex6Y5y8rVFwSol8LlTQ1My
CPzeTAFe5blhQqNL5rw82ak4B+ROn+a+n+ue6p+w22RmnejeWXaCOPg76b+FEicXim02M64nzEFk
cbNT1DPz/yE1RfoglvudVYgMvSv9mW0nvKxcn3r++MDv8wxB9FMWX9vF0XNzMob9nXN8pfZslJya
IYhaZFnEN1ruSce+PLqIf/AA9X91er/Wqqdy+SrZKrh2k8CKtgrWFzz7+Jze4ydFsjbYsnR+of6j
gMCRXg9wLzBJz2ULUNuMefN+c8PbMayWA/1SEBdXOsJaW+pKXwJAyadIo9tGTGd5DTnA+tYphB6h
9uYGCqse/6I90A+Nj63qVCoxJmD+rIrunC7G1c03umzPNxktcHao1dzU/BMvh31Y7f/ya7zJCO3u
lklbuJTCELlPiaAfLXiniwIavZE0ZnLqXRfUomHRxOJhzWJbAjk0xfa3w4oOdPtWM1JHE5r8bMMJ
CYQSKFEOMLbrh0IZJ7dv4eJBC/9D5me7HbS57/c2WNogqjDIa4TOy5HTHBTE/x9/rDvVsH2IIbac
chokQQ/f5Ghr2JMbfqT1ez41F1tMWwxw+v2YIi6H3TPgM2MXRQk4zrGADxtWu445v3WaPtLjKe6g
O4VFXGR8n9E/tqJ5EO53CeuaIOIRHSzJirpIdtbqTUNqXS60xezeah0i0jgT2xQ3h1Qn6hesV71P
gk4kyTdHqLS7RBD0qnVIxepAQtCkbxLV15JDMeetXmr5WHG0ekkEUTCXf66kkbZCT1v91adhqlaE
ws+JjggLdpKn+SSptLPBokmD+I7G/y/8DmcwPQYVZoKHhCPRjxLnEmEmcMU1MXisAicHIbCve8GO
/fC8/s1VboMGGXhi1sP6UwKB4/Qsi6d4ozZW5QFN+xLg0YeuXoaF9f8q4rbQdWEijcnaJQunxFGe
PtGyj96y1ebHT2/MBKne9eSDCGSCsAlXnAbd8t4uGOvJ8Kvsu8YiWyX+JO0f/FOp14xHI4yd8kSw
qU0g7u6p1zzndrZxeYBx96Bsmih01gBQQctwYpDkSK5HufQ/cKnBEkVp5JR1ZOwd2piTgrhT0nXq
3EeXnXjZ7pdCLrUSrJd75eun75tOj5rWtrps50hJsxHag4itaD9Jk37TQWaKXUuMucs8edg67St4
fRzTjFbU+rGUTSm9w3cXIGrCdNpGDSHMKpVdZT8YVBsIPjzBmN7vQ2NhGLlqzNZ2nloaCYCsOTVV
C+fofndhdaVFfxxr6CNDnl+0ppCvpCJPniACx37cqrH1uHu0eNzJSQfwKbBaZ+zEBYLc0LWg+YFm
hGfKjI8RXN3s4KpYWvDIbkODv/Yznl+GRu8MJJEV1SSurmiaBymlrqT6CLOxNHqyury60lCl7G46
ArG8wh/mQ2NLmZPOy/5n3hY9B+jaPwQAK56laR9T9p148DcpffGOWVT5v/bnj5mU6iybuRe+Zvz+
29SHxuKf97lVg5cetLLQTtLh7avyejxJROgsqV2nLJC4JKo+pAy95G9A7Im9cF37EWl2+a2dx0Mh
uiwrqqJyma4SbQyl4nHZVxNqHGLFXGLQB4UdAwdLWPn8nb3q8BbhVMuIBdagu+2ejvyCC5PfVYG9
4evEYIcWv37DVTsZTtAa5/cRJClCewie+z2HUYRjksd6DmIyuUWk/AuCZP6msRzsfhwfOz2rdPIt
G+TuChWUyHk+bURfXChWJwlUCNF8WDYcgqXyGGECUYLAfoOUyg4/32Lq+dPPBjLgsQR2xWAjQkvD
8uIsGu88ShbxKcfqhVrxpWVI13+NsogBSgxoJXUU/AYdSW9el3Ew3Ghuitvk6XpF86I9akNSS+nt
QBkd8Fb9GsPuG6JrZS2VIt6ev7CTVUfhTuRl33y1N+OnCznS8NQ+gW/37mi5LkNQLyIU9pCpeqpO
2P5aTywFSSsu1Z51cI+k4KWV3I5hH2WNueGDG4uWHjMlLeP8AGLmeOCu6kenX6a58oZZlrMlpktE
Cp5juzmMjuDii2B97mSirCrgfLWmfeIzpGhGqphXYRPEkYcOtSjWEHnLVQxNmkXDqM2D2it+24MM
0+wPomMSkpt2ZX4KineZ6AE0ziNnHKz/ewJEwUgnkHImDFnMYPgpISX0MgIBSb9Mrnyp5R/zPKId
ngjJzKrgRHGOLKq59SJWxdyeanssQf7sll+SVUuirHy0jTs1iEtALwsAl9mvBb1IQ4OT8r9yQxLh
UpBxVoqDirFWDRCe+sP0mLnxtU6vZnIIoND/HEqSqo566gRT4obAwXvvp4Prwh8m+LvJliJwGLdG
dVB3QjPkR2aSMdIy7WA9rmAuR8mrMHnORi8ULhTmtxAl8p4onW4rAkBfNPzXHoy+4x34cZJBGEU5
wnoiucalbcwip/x3cam+OjCRNDfxgXNyj7HpYQYwRTseKLyKjYAzdrAxyzQvbOgahnRbNtzIvMeD
MZG1BKdUQQZr+y08rF9akGGhYJviYJ4kboIAnrtz+rw8ucBBgEYeXo+wfYxBIzU9tt/V/RV1dtMZ
Ilg30D+aaImI7cxz/RXO4qa1PONU9FlUx3qOtTPeUOob7x/XNK1C+5g6YGIJZM2zey9DTKE2Dve0
GkG7ZZxDrU3AnGX2FRkYoywhVnMp6BwiT8cbL7Zd7U6dF65Sxi8wYtsram3VZ5k8IQH3yEpRLuLN
mV78S1fHM1fm/zv6sXzpr/Eu7C6/i89i9t1AwaeQNbDljrUA1YPXIpPwLgAgt4SLRBRAN+gTFcoF
+/8vVDogmPfd/0ghbH07/aM2siAKDpbWXH26MK62GGBzSxEmz5m5b5tahIYQELO3dXhBn9kY+W/g
JfrY9Be++WR9PsIZQTvxA75Bwp40eWBzBvbcxbslQytST5ajIS9TZ67RZ4p3jsRLTa3bZDAl5RC/
c1kXbE/KdIOKGTDFUxrqLrcsTom6miH7TD4744ZO4lYWxSP1q9LgXvEawH4nGF6fD6f0muIups1f
pdgw8jMNJDCteJBAE3MSwW7wqWnXI8ZrBlmdwk/GGtJTW8fH905LDrBJcHkjvyOwkcyhY240pzYQ
K1kYYOp7nIrNbJvIlIWzweJSTEIZhOLLJSZj7jLcKZeM7veEtsWlfw4+Ku1YJMj1e+OEa2kQw48u
+oQMH5P2HsPgxpgVdAjjnOYTzWvRvLjbZsH4So3F4G9W
`pragma protect end_protected
