`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
JFT7olhrsTCn+ua1lge2xzJc6xV9zehjCT5vMCN6GPUIf8dvvCgCGnH0PryzpF2T3u8VgDN2GJ1d
OEw+xSU4XQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DWN4fzIO1W1DFLPBoYl4OYwBRXztzK+LBLr4z1/82R1MFFbfQvskKIvCWAR1MRziyWgaYO9LnzdX
xA7PpBQLU0K79QvubOk6+a1Ss5+eO9Ildkm7dEXBb9XwHNBHUMhEH1bMJRHMA7tfx570l4MEM/yL
5BJy8k1v9ZEb1wyr7fw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
GsloE+YSC8eF8ZjGMHJ9cowlE4zZtchVLe39wyJxfV/9Su4KfXPknTKrqPtB7w75vtJ6aUF5WgsZ
D9WzwYFAkocFRmoBZGcZpl9cKg1+oj2xsKxv4CyJjZrIfriVNBoQsjv3mv2Pl1cUU6whc+VGaZ2S
WQqq0AGeen3e5hh2jR8C6VcXmzNUEOpUXGJXdLs8uTMLVNhDrRGT52GKlJwAauElnA1GRZlDU/4P
tduimEh1lJxNW9cQKrEhyaw6GHOKSpCQYKa6iz2hcaTTM5ukIifpRBsViA9EA019NKau7wX5do15
44WrGQ6Pku2+p41P5gXXGoIC9PJUqOVHrJJqvA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dm2h0SfQUU6hjNgoA0pqw4ElcOLURiRQMlNp8Ljva1cvpbZdr23LtP2d8w5NNgrg4ofcEkTfPoCi
qeFAQgrfNAYSAHzgC4BJaxJwYs9imY4ko6Sy1O42y0az8iGpGoKBSvNSX5xuLUjwPt785DF7bxnT
pJe3l4kU/rKQ/JHJSYZDavZhz7Lto2otnDfEKCpKOHR59wSuCDIJFV9vgrCQJiMLGTLRYl+Q057D
cARSN+sOdWxzBHZdChGlYm9NS44xOvOnNqQPykmp87UohNE5kXrEfABQHVlCHBrp1yNnZwGPmB/0
EWp+59x7lh8LJKJv2R+xoENeBLJSbODhJrg+zA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KLXlplMxMOr1UBh/V5AsV69JA8GA3+Vp5E8rfDFcFwrKpB0qUC98FVfyYjX0wZ7hvcN0+jIU4kWT
vFIuyoldYnLu7XbvYamToCH9VsQSxHreBi3oMuK7rcmOPb4y7t0YHitun763RL73Fm9GWd2IEjlU
HOmVreB8GHjZEMSCjh6O39X0h4Xb4LfoWf0i6Bg08GyZ3e+Rbvu4NPstL9O+YLzBTo2FvlWx9JZU
7OWmMADvdgLxnJDZC7hGmOW1pFgsEVLQYNOnmSPpBLU7R/oDo12I2dfWTARjOaDdAGCKyXLK5uFD
b9957h/Z204aRFv25nyrJMZ0U0DgVcbsJFjaeg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
i8S77Q8PhqhUkfeFveat2i35TbsLYBPdAL2QEQ24FrUhgbaJI98QdPzn95fQYWjX8bBYO6c7S4gI
XiyWHFsxrYW9TGaKwZYZ2HLQIYrp+WDKsCsXA/CidvbAZW+M2UelTLU+isKkz7R5gdwrMiFTa6/J
LJf6mpx/GKxxwOfMNnc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Gu0KbdM1rFg2ntk8q9kyOlc0bktBZ3dwHmgv3XVJwWJJ/JvhU1/FpUsRHKoW3jrRV3KqhkKbHHap
qmHQ3yAa5guKP9HWchAtStr/o/5/gykqC/E9gv5nOb9WTzVEnIuivDNYb3V1jYeiUwp1D1udgk1c
e/UQbOJ1prqLDgwjmJHJnbgc6vStOjj4AwjvAnAYPJiolFJIVScEp7Lk7zWE5wY164tJV7VT3hPV
GG5rJM3+KZUD8K1NQfH3EpQsi2yar+87kFlgJznKw8ABh/jZe5skBIXFxZOHuK0ihGEH/KNJ1wVl
2WA2hx5dSaQuxCSLW3A8LUpsdcC5JHh16ITaNQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
/uyJlef/Ij1AWiQn0ynjAcNR4xRu6tMAHifLxAVQEI+G9yNscU8+3BBvfZXI6L0PkAPvv6uiQUPZ
DuGYHN/e/S9IgxrXjSzp/lYlFPyXCsxAcTR26wqTzqsZ4EjPB9ffs+666dZqZds1Zk4DkYFvIyhy
3p0YtKjVFYNeRQAzlWupPlaSHP9VurkwU7JSeeshjbhvDg8UgcL1idSWEzEuIlaE8ok7y7Sy5U4F
uqxYo/kiALBMq6yf9RCUyH+GtgQDIXnUHyauHSUythXF7K5SQSdokLvihpm6lKhVKYnT9lAqHHis
PV7Bv/kE1RBrtp+nJJryDNfU7gvJ/TMlu06SbjLADNoCeN+oI/B3z1cGL6lKYhplpd+uhkwno9E/
MP9bFnzEpfckmgjVGXkSnsDUOTxuZsfGjtzukHYvzm40opNyAh4M2ZU0rzWfQkJZ5FGqqJogUwiV
8Pio/ouU9JBE+KvCpsojtf/uQNwjJluHleoE68IX1LdsJLHm2e9hK3esDwBkxdyNc7BafCoRzNrX
2KczzIN8XvH9BMz4DTdZT07XvgJFz+GrfuDkl+sVSUGfzZrCsvsx1gmfaytxz6BUv7qJI5DN+8RR
FXXZjyczq4XJKIicRiHle8qi5mizahMBeijXD1DxyKELbOCrbrVTSB98iP5mU/fElI7SFFpLWvU3
x4ZjizTD7FjGJAiein6oxY+DBNAnTpTIRXjsnP4mTPrmSV32EpCp/0bMY1OS7BYsM0QvsOcCZoAH
nVK1X/LSdoq70A7/J1UkxsZ6zqK2Bb5UCTTn/n/Dmy+EqsooRzc+QZCDnnQogzLsQ+YcVEwn7fRj
6YvoLcuSRwpo/oBkyg5BB+mzR1XLLjSK8rgf3WZIrIbCv9qeTH5G95MVqRG+P83nxFKenZACf5uv
5DZW/+T02FFs19ab+2D3WckGCwKctTms3W6bGMR6ywQGCcc5mWMMwlOHHI7uNMV/L4jad+9BrJ1E
hgsq4bS28zEFK7yWffd/zS0q3ZuS82ekjZH0MnNN7cuzammQtjYUgO0A41ftEo0K0llaWj4jiBYb
MDYQVc0weMLG+mv4kDKiUijQshH+94DKdYVqOyVbuFjYxrTXmwlLavWgsd6cngAzAmuZ4G9EmGWz
QCA8DHlPfUMNExZCYoRtGH5s3Feaw7k2ACIjydh05RnXyuPx7iYBl19cinhwlYlIg7Sqk9F6qpVd
IBgvI6Z9s5/e2uIZUj+QY57OAEA0LKBgRYNsh/dLGHm4y4VvqAACy8UbHGKKrokGYwWb9C+vnM9x
cfm13eGiV2YXdM4SiGF7tbPrmJ2hxFj1yq2s28FteJfW2pSug3NXgVPv0MF++AplLP2feFLqqqZa
fFE9APU+Qp2bIl32NL16Nt4EX75OhRs19mZpn4xiXvkH4z4XfzkP4CeuEc4qZHSjWz+gQMkuesjV
LD3Az7UEwW76BcsycoMH1rFREaoHtfVjEQ1OaaGXRXXyaavtEOQG5ptIrffe6kKfWFc1Sh05vBJQ
YvbwZIsyZ+3a3j53OgIAdWAVsZiTDUI1+vsGuRhIreL/FY7Ry8ahw8aZn7ky5rvUbiH10CC+TXRT
aPV1m+dDb1NnoELmtf6PIjElz16tRGb5RnEmOxeMklvfveuyXaRsTionxLpKvLx6EmaHQI5Q1W95
lRRp5CtrSavp2tDa/c+DZWvLx0i2HyBNxcUx/OEOvFxaN4q/ufgOxHI+rhBzMJNrTAr32H5g/USe
S4G+MdHpZnxtZyghtCsMDGGkmtnnJbpNW3DCuyDHEsSncZik2fnOu1i1BTC7wyr39QOo6udhsc1d
j+Nl20EX7PXJA3iijEiibJKjcVud3KhrZFNdMCmGBi0ClO7uyCaOfm3GhZojpVqs3V1mHFJb1xWI
j/bk+wXaEFIN7TGMCn1NG57JiJhD6P+fNzJQDPl2YY04CSJEy12bigWmSFZHWqPWzpdSJ6a1Vpez
9ZJCC0UDZq5xVBfW5s1B1G/j3CzbHbt3LZ6ss4pK+ffPECFmsLmuGbKEA6/7908W9fnWqTrAP43A
CerePBJ3pyN1GXI1cVRv/FEQbnynESTBQDhmYencDv9jcn1rOsTOz1w/u4CIAvcWb3Ohi+2tSVz6
v365I0+5a44KoQcyxxNL8JFxCK2bAtxqZsVdtbpci1RDJJbXBKE7fr92SFzIeJDho1LH4OGUUFUo
34B0KYc/knSoTQaCP5eEqIkLaqJIwI/U1Zy5sbwftub1N8OPzxUwG7HH9W2LxymNXuf912e325J1
OgNAGX0at6AIfeAxWiAPfGrvUs+pfSVMeu/L/hYxpzNCV43xtnkwJXJWXRQ7LNJ9DpSkrfGzOuNp
AEeW0AGXQaHUMPKqoVYZKUnxDDxDrrtJQJeiWrYXl9XVZir1nwxJwqWtRHN+TrfOSTMJkPMojO7G
ppb9hPTDDC0/4MRmvh74ee+Q9o8RrZjiwU86xkjw9aVk8OAwrm3YqLexwFo7xy25KwKi8SJeDKrm
xa59qeltNpIDb+oo1KllIoV7kE+QrOPXatdYa0Mk2Br2ENSSCkrrtyweMvHrmh577iUUHHn1hYba
AAJyXApzpc5Zj8xjkropP9AhbIJ0Ds1mVJh9VZEYVHu6MOuZOP4jeBfUwnvkprUPB/nyDYT0wX3J
O0fp9+TYIUC/LnYFhMskK7wur17Tes7e/ZK/JrMPzgua8ak25cx22J8odHpiQczsPH/0ed16TVsO
069zyKCsdhWl4ZkPhUrZWlE1cLsQtEG4TigOLHFXQzGtrUI52IgmfvS8amilXROaDkXNZH8gtUZL
DBmIUH++ISeoab5EZu9kucGGU0qtnirPdqMx1iaJkA2W0bhrQM9L5yvSBRGnoI5jkiZSQxCs2Jad
RXxRlaMbO0lWoW+NHLenmlCZgg8kdtizLBwakmObmFMEftOucUeB4VpM/UjeM14iiYAUyfhooxzA
CwSXs8DS3UBL1THmyCgUxVaTVCQzZ4NuOkDodtO9U7tGib0NrsHp1IItrdS3aYZ2xIASoEBJKuCA
/vgbd48vkNy7FZ6m/xENerJgaguQZFEUcWcQrabVh5DhNKCYkuHVOcYFPGZMqNi8q49IfLghc58M
SQ0zoSSecM8RlU+eyx3MKvAtLJUievVGDyj2Yx3aJlTrGlMaETAjj4RM9ZNiwpcHeHXZtYxS80Ri
IOKgrDXHf5ATWvM+VPNtlXTXAQV0rH9rA3q3ankXk/qYsPSpGZJdTqY/rNVg5H6YacKrJyswMW5E
0eZ72eEduNdhLMWFzpnflKR9J9FccF8xS56URIRlhGQjG+KnvRiyfLS+RIVa5VJziuGQSbFLAnKk
1s0QjywE4mKmS0xr4qfYqEpUQJcd54urK2XU05JfOS0qx56llE4oEhmKTuaQU4D9CqClR5zjwZ2I
sbld9J7JLHOSxyPifDqd9BB+DW6i4R3nQ+sY46LFMWD3kvSUkNLi3Y+JjWudmC2npwrrHTV/4Xcr
ZPL+dl8tY6qaGWbZRHMNPdJM4QFO/vyx5v0zDNFteaVhNUynKoQGWafczZEO4abyO6dDgQ6bKv+H
AopJLcmauGaRyuyxAdlskPeTlJCY2Ics71I7sD6WS9xhome58G1aOfagNUkxTknGIQS+IWlzOjol
8ihDz+S9elJNltQCBZA5N670l9/5QUxoOtyBrRSUC1z0AvfFBlwp15tQhI9NpniMXdZfDVvBBBtU
8dAkX00NfHdyBd9+VY6PBnHvKAiOtrG1BJVFaILINRWPnSRkApAbjhve+zGUd2+pEYayQu099L1E
1WYZRKPEqYmOdUbpzWMqEyb18bNYdzauoVEnuMobzyVEB1UBfQ5GGRt/FDbTAjSkLsay8lrST79V
TzQJCREBl1DAUbZJW3IWTYNN2Muj+V9XSztqcBDaxoIouAPwXEGPye01UivI8yKmMa1OqmaJdDaP
F1zhW3wJq1k5d1tRTxLWjKMos5t5Ui1Q7/uXiNnbCA0dJq8B65fwxOUGZu16etGWT6XAmwKlb+pZ
SjW8xb6WVqemu7dAOvdZnhW+gQKTcDTqHRooP04IJ9wNuEEqEK2eA/pg7HvQ+2TYnqdtvMBFnF+y
m+XimV+RFyroRQ4EStBgm7RTuyiKSsNKF599YZDlOvikFCUo31YLzVtg8HZEssv4Nc4T7oRQj6Gg
kg==
`pragma protect end_protected
